magic
tech ihp-sg13g2
magscale 1 2
timestamp 1766118055
<< metal1 >>
rect 1152 12872 11424 12896
rect 1152 12832 3688 12872
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 4056 12832 11424 12872
rect 1152 12808 11424 12832
rect 2851 12536 2909 12537
rect 2851 12496 2860 12536
rect 2900 12496 2909 12536
rect 2851 12495 2909 12496
rect 7459 12536 7517 12537
rect 7459 12496 7468 12536
rect 7508 12496 7517 12536
rect 7459 12495 7517 12496
rect 3235 12452 3293 12453
rect 3235 12412 3244 12452
rect 3284 12412 3293 12452
rect 3235 12411 3293 12412
rect 3619 12452 3677 12453
rect 3619 12412 3628 12452
rect 3668 12412 3677 12452
rect 3619 12411 3677 12412
rect 4675 12452 4733 12453
rect 4675 12412 4684 12452
rect 4724 12412 4733 12452
rect 4675 12411 4733 12412
rect 4875 12452 4917 12461
rect 4875 12412 4876 12452
rect 4916 12412 4917 12452
rect 4875 12403 4917 12412
rect 5059 12452 5117 12453
rect 5059 12412 5068 12452
rect 5108 12412 5117 12452
rect 5059 12411 5117 12412
rect 5355 12452 5397 12461
rect 5355 12412 5356 12452
rect 5396 12412 5397 12452
rect 5355 12403 5397 12412
rect 6019 12452 6077 12453
rect 6019 12412 6028 12452
rect 6068 12412 6077 12452
rect 6019 12411 6077 12412
rect 6307 12452 6365 12453
rect 6307 12412 6316 12452
rect 6356 12412 6365 12452
rect 6307 12411 6365 12412
rect 8707 12452 8765 12453
rect 8707 12412 8716 12452
rect 8756 12412 8765 12452
rect 8707 12411 8765 12412
rect 4971 12368 5013 12377
rect 4971 12328 4972 12368
rect 5012 12328 5013 12368
rect 4971 12319 5013 12328
rect 3051 12284 3093 12293
rect 3051 12244 3052 12284
rect 3092 12244 3093 12284
rect 3051 12235 3093 12244
rect 3723 12284 3765 12293
rect 3723 12244 3724 12284
rect 3764 12244 3765 12284
rect 3723 12235 3765 12244
rect 4003 12284 4061 12285
rect 4003 12244 4012 12284
rect 4052 12244 4061 12284
rect 4003 12243 4061 12244
rect 6411 12284 6453 12293
rect 6411 12244 6412 12284
rect 6452 12244 6453 12284
rect 6411 12235 6453 12244
rect 7275 12284 7317 12293
rect 7275 12244 7276 12284
rect 7316 12244 7317 12284
rect 7275 12235 7317 12244
rect 9379 12284 9437 12285
rect 9379 12244 9388 12284
rect 9428 12244 9437 12284
rect 9379 12243 9437 12244
rect 1152 12116 11424 12140
rect 1152 12076 4928 12116
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 5296 12076 11424 12116
rect 1152 12052 11424 12076
rect 1899 11948 1941 11957
rect 1899 11908 1900 11948
rect 1940 11908 1941 11948
rect 1899 11899 1941 11908
rect 5923 11948 5981 11949
rect 5923 11908 5932 11948
rect 5972 11908 5981 11948
rect 5923 11907 5981 11908
rect 8515 11948 8573 11949
rect 8515 11908 8524 11948
rect 8564 11908 8573 11948
rect 8515 11907 8573 11908
rect 3531 11864 3573 11873
rect 3531 11824 3532 11864
rect 3572 11824 3573 11864
rect 3531 11815 3573 11824
rect 1219 11780 1277 11781
rect 1219 11740 1228 11780
rect 1268 11740 1277 11780
rect 1219 11739 1277 11740
rect 1411 11780 1469 11781
rect 1411 11740 1420 11780
rect 1460 11740 1469 11780
rect 1411 11739 1469 11740
rect 2179 11780 2237 11781
rect 2179 11740 2188 11780
rect 2228 11740 2237 11780
rect 2179 11739 2237 11740
rect 2851 11780 2909 11781
rect 2851 11740 2860 11780
rect 2900 11740 2909 11780
rect 2851 11739 2909 11740
rect 3147 11780 3189 11789
rect 3147 11740 3148 11780
rect 3188 11740 3189 11780
rect 3147 11731 3189 11740
rect 3339 11780 3381 11789
rect 3339 11740 3340 11780
rect 3380 11740 3381 11780
rect 3339 11731 3381 11740
rect 3907 11780 3965 11781
rect 3907 11740 3916 11780
rect 3956 11740 3965 11780
rect 3907 11739 3965 11740
rect 4771 11780 4829 11781
rect 4771 11740 4780 11780
rect 4820 11740 4829 11780
rect 4771 11739 4829 11740
rect 6123 11780 6165 11789
rect 6123 11740 6124 11780
rect 6164 11740 6165 11780
rect 6123 11731 6165 11740
rect 6499 11780 6557 11781
rect 6499 11740 6508 11780
rect 6548 11740 6557 11780
rect 6499 11739 6557 11740
rect 7363 11780 7421 11781
rect 7363 11740 7372 11780
rect 7412 11740 7421 11780
rect 7363 11739 7421 11740
rect 9379 11780 9437 11781
rect 9379 11740 9388 11780
rect 9428 11740 9437 11780
rect 9379 11739 9437 11740
rect 9579 11780 9621 11789
rect 9579 11740 9580 11780
rect 9620 11740 9621 11780
rect 9579 11731 9621 11740
rect 9763 11780 9821 11781
rect 9763 11740 9772 11780
rect 9812 11740 9821 11780
rect 9763 11739 9821 11740
rect 10627 11780 10685 11781
rect 10627 11740 10636 11780
rect 10676 11740 10685 11780
rect 10627 11739 10685 11740
rect 1699 11696 1757 11697
rect 1699 11656 1708 11696
rect 1748 11656 1757 11696
rect 1699 11655 1757 11656
rect 2955 11696 2997 11705
rect 2955 11656 2956 11696
rect 2996 11656 2997 11696
rect 2955 11647 2997 11656
rect 9675 11612 9717 11621
rect 9675 11572 9676 11612
rect 9716 11572 9717 11612
rect 9675 11563 9717 11572
rect 2091 11528 2133 11537
rect 2091 11488 2092 11528
rect 2132 11488 2133 11528
rect 2091 11479 2133 11488
rect 3339 11528 3381 11537
rect 3339 11488 3340 11528
rect 3380 11488 3381 11528
rect 3339 11479 3381 11488
rect 8707 11528 8765 11529
rect 8707 11488 8716 11528
rect 8756 11488 8765 11528
rect 8707 11487 8765 11488
rect 9955 11528 10013 11529
rect 9955 11488 9964 11528
rect 10004 11488 10013 11528
rect 9955 11487 10013 11488
rect 1152 11360 11424 11384
rect 1152 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 11424 11360
rect 1152 11296 11424 11320
rect 11107 11192 11165 11193
rect 11107 11152 11116 11192
rect 11156 11152 11165 11192
rect 11107 11151 11165 11152
rect 5827 11024 5885 11025
rect 5827 10984 5836 11024
rect 5876 10984 5885 11024
rect 5827 10983 5885 10984
rect 1987 10940 2045 10941
rect 1987 10900 1996 10940
rect 2036 10900 2045 10940
rect 1987 10899 2045 10900
rect 2851 10940 2909 10941
rect 2851 10900 2860 10940
rect 2900 10900 2909 10940
rect 2851 10899 2909 10900
rect 4387 10940 4445 10941
rect 4387 10900 4396 10940
rect 4436 10900 4445 10940
rect 4387 10899 4445 10900
rect 5451 10940 5493 10949
rect 5451 10900 5452 10940
rect 5492 10900 5493 10940
rect 5451 10891 5493 10900
rect 5539 10940 5597 10941
rect 5539 10900 5548 10940
rect 5588 10900 5597 10940
rect 5539 10899 5597 10900
rect 6403 10940 6461 10941
rect 6403 10900 6412 10940
rect 6452 10900 6461 10940
rect 6403 10899 6461 10900
rect 7563 10940 7605 10949
rect 7563 10900 7564 10940
rect 7604 10900 7605 10940
rect 7563 10891 7605 10900
rect 7755 10940 7797 10949
rect 7755 10900 7756 10940
rect 7796 10900 7797 10940
rect 7755 10891 7797 10900
rect 8227 10940 8285 10941
rect 8227 10900 8236 10940
rect 8276 10900 8285 10940
rect 8227 10899 8285 10900
rect 8515 10940 8573 10941
rect 8515 10900 8524 10940
rect 8564 10900 8573 10940
rect 8515 10899 8573 10900
rect 9091 10940 9149 10941
rect 9091 10900 9100 10940
rect 9140 10900 9149 10940
rect 9091 10899 9149 10900
rect 9955 10940 10013 10941
rect 9955 10900 9964 10940
rect 10004 10900 10013 10940
rect 9955 10899 10013 10900
rect 1611 10856 1653 10865
rect 1611 10816 1612 10856
rect 1652 10816 1653 10856
rect 1611 10807 1653 10816
rect 8715 10856 8757 10865
rect 8715 10816 8716 10856
rect 8756 10816 8757 10856
rect 8715 10807 8757 10816
rect 4003 10772 4061 10773
rect 4003 10732 4012 10772
rect 4052 10732 4061 10772
rect 4003 10731 4061 10732
rect 5059 10772 5117 10773
rect 5059 10732 5068 10772
rect 5108 10732 5117 10772
rect 5059 10731 5117 10732
rect 6891 10772 6933 10781
rect 6891 10732 6892 10772
rect 6932 10732 6933 10772
rect 6891 10723 6933 10732
rect 7659 10772 7701 10781
rect 7659 10732 7660 10772
rect 7700 10732 7701 10772
rect 7659 10723 7701 10732
rect 8043 10772 8085 10781
rect 8043 10732 8044 10772
rect 8084 10732 8085 10772
rect 8043 10723 8085 10732
rect 1152 10604 11424 10628
rect 1152 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 11424 10604
rect 1152 10540 11424 10564
rect 1323 10436 1365 10445
rect 1323 10396 1324 10436
rect 1364 10396 1365 10436
rect 1323 10387 1365 10396
rect 3435 10436 3477 10445
rect 3435 10396 3436 10436
rect 3476 10396 3477 10436
rect 3435 10387 3477 10396
rect 4867 10436 4925 10437
rect 4867 10396 4876 10436
rect 4916 10396 4925 10436
rect 4867 10395 4925 10396
rect 5059 10436 5117 10437
rect 5059 10396 5068 10436
rect 5108 10396 5117 10436
rect 5059 10395 5117 10396
rect 5827 10436 5885 10437
rect 5827 10396 5836 10436
rect 5876 10396 5885 10436
rect 5827 10395 5885 10396
rect 8803 10436 8861 10437
rect 8803 10396 8812 10436
rect 8852 10396 8861 10436
rect 8803 10395 8861 10396
rect 9955 10352 10013 10353
rect 9955 10312 9964 10352
rect 10004 10312 10013 10352
rect 9955 10311 10013 10312
rect 1507 10268 1565 10269
rect 1507 10228 1516 10268
rect 1556 10228 1565 10268
rect 1507 10227 1565 10228
rect 1603 10268 1661 10269
rect 1603 10228 1612 10268
rect 1652 10228 1661 10268
rect 1603 10227 1661 10228
rect 2755 10268 2813 10269
rect 2755 10228 2764 10268
rect 2804 10228 2813 10268
rect 2755 10227 2813 10228
rect 2947 10268 3005 10269
rect 2947 10228 2956 10268
rect 2996 10228 3005 10268
rect 2947 10227 3005 10228
rect 3907 10268 3965 10269
rect 3907 10228 3916 10268
rect 3956 10228 3965 10268
rect 3907 10227 3965 10228
rect 4195 10268 4253 10269
rect 4195 10228 4204 10268
rect 4244 10228 4253 10268
rect 4195 10227 4253 10228
rect 5163 10268 5205 10277
rect 5163 10228 5164 10268
rect 5204 10228 5205 10268
rect 5163 10219 5205 10228
rect 5259 10268 5301 10277
rect 5259 10228 5260 10268
rect 5300 10228 5301 10268
rect 5259 10219 5301 10228
rect 5355 10268 5397 10277
rect 5355 10228 5356 10268
rect 5396 10228 5397 10268
rect 5355 10219 5397 10228
rect 5547 10268 5589 10277
rect 5547 10228 5548 10268
rect 5588 10228 5589 10268
rect 5547 10219 5589 10228
rect 5643 10268 5685 10277
rect 5643 10228 5644 10268
rect 5684 10228 5685 10268
rect 5643 10219 5685 10228
rect 5739 10268 5781 10277
rect 5739 10228 5740 10268
rect 5780 10228 5781 10268
rect 5739 10219 5781 10228
rect 6115 10268 6173 10269
rect 6115 10228 6124 10268
rect 6164 10228 6173 10268
rect 6115 10227 6173 10228
rect 6979 10268 7037 10269
rect 6979 10228 6988 10268
rect 7028 10228 7037 10268
rect 6979 10227 7037 10228
rect 7179 10268 7221 10277
rect 7179 10228 7180 10268
rect 7220 10228 7221 10268
rect 7179 10219 7221 10228
rect 7651 10268 7709 10269
rect 7651 10228 7660 10268
rect 7700 10228 7709 10268
rect 7651 10227 7709 10228
rect 7747 10268 7805 10269
rect 7747 10228 7756 10268
rect 7796 10228 7805 10268
rect 7747 10227 7805 10228
rect 8131 10268 8189 10269
rect 8131 10228 8140 10268
rect 8180 10228 8189 10268
rect 8131 10227 8189 10228
rect 9195 10268 9237 10277
rect 9195 10228 9196 10268
rect 9236 10228 9237 10268
rect 9195 10219 9237 10228
rect 10243 10268 10301 10269
rect 10243 10228 10252 10268
rect 10292 10228 10301 10268
rect 10243 10227 10301 10228
rect 10443 10268 10485 10277
rect 10443 10228 10444 10268
rect 10484 10228 10485 10268
rect 10443 10219 10485 10228
rect 11299 10268 11357 10269
rect 11299 10228 11308 10268
rect 11348 10228 11357 10268
rect 11299 10227 11357 10228
rect 7083 10184 7125 10193
rect 7083 10144 7084 10184
rect 7124 10144 7125 10184
rect 7083 10135 7125 10144
rect 7939 10184 7997 10185
rect 7939 10144 7948 10184
rect 7988 10144 7997 10184
rect 7939 10143 7997 10144
rect 2083 10100 2141 10101
rect 2083 10060 2092 10100
rect 2132 10060 2141 10100
rect 2083 10059 2141 10060
rect 9387 10100 9429 10109
rect 9387 10060 9388 10100
rect 9428 10060 9429 10100
rect 9387 10051 9429 10060
rect 10627 10100 10685 10101
rect 10627 10060 10636 10100
rect 10676 10060 10685 10100
rect 10627 10059 10685 10060
rect 6027 10016 6069 10025
rect 6027 9976 6028 10016
rect 6068 9976 6069 10016
rect 6027 9967 6069 9976
rect 9771 10016 9813 10025
rect 9771 9976 9772 10016
rect 9812 9976 9813 10016
rect 9771 9967 9813 9976
rect 10347 10016 10389 10025
rect 10347 9976 10348 10016
rect 10388 9976 10389 10016
rect 10347 9967 10389 9976
rect 1152 9848 11424 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 11424 9848
rect 1152 9784 11424 9808
rect 4003 9680 4061 9681
rect 4003 9640 4012 9680
rect 4052 9640 4061 9680
rect 4003 9639 4061 9640
rect 4395 9680 4437 9689
rect 4395 9640 4396 9680
rect 4436 9640 4437 9680
rect 4395 9631 4437 9640
rect 11011 9680 11069 9681
rect 11011 9640 11020 9680
rect 11060 9640 11069 9680
rect 11011 9639 11069 9640
rect 1219 9512 1277 9513
rect 1219 9472 1228 9512
rect 1268 9472 1277 9512
rect 1219 9471 1277 9472
rect 1987 9428 2045 9429
rect 1987 9388 1996 9428
rect 2036 9388 2045 9428
rect 1987 9387 2045 9388
rect 2851 9428 2909 9429
rect 2851 9388 2860 9428
rect 2900 9388 2909 9428
rect 2851 9387 2909 9388
rect 4299 9428 4341 9437
rect 4299 9388 4300 9428
rect 4340 9388 4341 9428
rect 4299 9379 4341 9388
rect 4483 9428 4541 9429
rect 4483 9388 4492 9428
rect 4532 9388 4541 9428
rect 4483 9387 4541 9388
rect 4675 9428 4733 9429
rect 4675 9388 4684 9428
rect 4724 9388 4733 9428
rect 4675 9387 4733 9388
rect 5059 9428 5117 9429
rect 5059 9388 5068 9428
rect 5108 9388 5117 9428
rect 5059 9387 5117 9388
rect 6211 9428 6269 9429
rect 6211 9388 6220 9428
rect 6260 9388 6269 9428
rect 6211 9387 6269 9388
rect 6403 9428 6461 9429
rect 6403 9388 6412 9428
rect 6452 9388 6461 9428
rect 6403 9387 6461 9388
rect 6603 9428 6645 9437
rect 6603 9388 6604 9428
rect 6644 9388 6645 9428
rect 6603 9379 6645 9388
rect 6795 9428 6837 9437
rect 6795 9388 6796 9428
rect 6836 9388 6837 9428
rect 6795 9379 6837 9388
rect 7459 9428 7517 9429
rect 7459 9388 7468 9428
rect 7508 9388 7517 9428
rect 7459 9387 7517 9388
rect 7843 9428 7901 9429
rect 7843 9388 7852 9428
rect 7892 9388 7901 9428
rect 7843 9387 7901 9388
rect 8139 9428 8181 9437
rect 8139 9388 8140 9428
rect 8180 9388 8181 9428
rect 8139 9379 8181 9388
rect 8235 9428 8277 9437
rect 8235 9388 8236 9428
rect 8276 9388 8277 9428
rect 8235 9379 8277 9388
rect 8331 9428 8373 9437
rect 8331 9388 8332 9428
rect 8372 9388 8373 9428
rect 8331 9379 8373 9388
rect 8427 9428 8469 9437
rect 8427 9388 8428 9428
rect 8468 9388 8469 9428
rect 8427 9379 8469 9388
rect 8619 9428 8661 9437
rect 8619 9388 8620 9428
rect 8660 9388 8661 9428
rect 8619 9379 8661 9388
rect 8995 9428 9053 9429
rect 8995 9388 9004 9428
rect 9044 9388 9053 9428
rect 8995 9387 9053 9388
rect 9859 9428 9917 9429
rect 9859 9388 9868 9428
rect 9908 9388 9917 9428
rect 9859 9387 9917 9388
rect 1611 9344 1653 9353
rect 1611 9304 1612 9344
rect 1652 9304 1653 9344
rect 1611 9295 1653 9304
rect 6507 9344 6549 9353
rect 6507 9304 6508 9344
rect 6548 9304 6549 9344
rect 6507 9295 6549 9304
rect 1419 9260 1461 9269
rect 1419 9220 1420 9260
rect 1460 9220 1461 9260
rect 1419 9211 1461 9220
rect 5163 9260 5205 9269
rect 5163 9220 5164 9260
rect 5204 9220 5205 9260
rect 5163 9211 5205 9220
rect 5539 9260 5597 9261
rect 5539 9220 5548 9260
rect 5588 9220 5597 9260
rect 5539 9219 5597 9220
rect 7947 9260 7989 9269
rect 7947 9220 7948 9260
rect 7988 9220 7989 9260
rect 7947 9211 7989 9220
rect 11011 9260 11069 9261
rect 11011 9220 11020 9260
rect 11060 9220 11069 9260
rect 11011 9219 11069 9220
rect 1152 9092 11424 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 11424 9092
rect 1152 9028 11424 9052
rect 1987 8924 2045 8925
rect 1987 8884 1996 8924
rect 2036 8884 2045 8924
rect 1987 8883 2045 8884
rect 5251 8924 5309 8925
rect 5251 8884 5260 8924
rect 5300 8884 5309 8924
rect 5251 8883 5309 8884
rect 2859 8840 2901 8849
rect 2859 8800 2860 8840
rect 2900 8800 2901 8840
rect 2859 8791 2901 8800
rect 3243 8840 3285 8849
rect 3243 8800 3244 8840
rect 3284 8800 3285 8840
rect 3243 8791 3285 8800
rect 3619 8840 3677 8841
rect 3619 8800 3628 8840
rect 3668 8800 3677 8840
rect 3619 8799 3677 8800
rect 5451 8840 5493 8849
rect 5451 8800 5452 8840
rect 5492 8800 5493 8840
rect 5451 8791 5493 8800
rect 8619 8840 8661 8849
rect 8619 8800 8620 8840
rect 8660 8800 8661 8840
rect 8619 8791 8661 8800
rect 11115 8840 11157 8849
rect 11115 8800 11116 8840
rect 11156 8800 11157 8840
rect 11115 8791 11157 8800
rect 1699 8756 1757 8757
rect 1699 8716 1708 8756
rect 1748 8716 1757 8756
rect 1699 8715 1757 8716
rect 1803 8756 1845 8765
rect 1803 8716 1804 8756
rect 1844 8716 1845 8756
rect 1803 8707 1845 8716
rect 2187 8756 2229 8765
rect 2187 8716 2188 8756
rect 2228 8716 2229 8756
rect 2187 8707 2229 8716
rect 2283 8756 2325 8765
rect 2283 8716 2284 8756
rect 2324 8716 2325 8756
rect 2283 8707 2325 8716
rect 2763 8756 2805 8765
rect 2763 8716 2764 8756
rect 2804 8716 2805 8756
rect 2763 8707 2805 8716
rect 2947 8756 3005 8757
rect 2947 8716 2956 8756
rect 2996 8716 3005 8756
rect 2947 8715 3005 8716
rect 3147 8756 3189 8765
rect 3147 8716 3148 8756
rect 3188 8716 3189 8756
rect 3147 8707 3189 8716
rect 3339 8756 3381 8765
rect 3339 8716 3340 8756
rect 3380 8716 3381 8756
rect 3339 8707 3381 8716
rect 3811 8756 3869 8757
rect 3811 8716 3820 8756
rect 3860 8716 3869 8756
rect 3811 8715 3869 8716
rect 4099 8756 4157 8757
rect 4099 8716 4108 8756
rect 4148 8716 4157 8756
rect 4099 8715 4157 8716
rect 4291 8756 4349 8757
rect 4291 8716 4300 8756
rect 4340 8716 4349 8756
rect 4291 8715 4349 8716
rect 4579 8756 4637 8757
rect 4579 8716 4588 8756
rect 4628 8716 4637 8756
rect 4579 8715 4637 8716
rect 5827 8756 5885 8757
rect 5827 8716 5836 8756
rect 5876 8716 5885 8756
rect 5827 8715 5885 8716
rect 6691 8756 6749 8757
rect 6691 8716 6700 8756
rect 6740 8716 6749 8756
rect 6691 8715 6749 8716
rect 8227 8756 8285 8757
rect 8227 8716 8236 8756
rect 8276 8716 8285 8756
rect 8227 8715 8285 8716
rect 8515 8756 8573 8757
rect 8515 8716 8524 8756
rect 8564 8716 8573 8756
rect 8515 8715 8573 8716
rect 8811 8756 8853 8765
rect 8811 8716 8812 8756
rect 8852 8716 8853 8756
rect 8811 8707 8853 8716
rect 8907 8756 8949 8765
rect 8907 8716 8908 8756
rect 8948 8716 8949 8756
rect 8907 8707 8949 8716
rect 9003 8756 9045 8765
rect 9003 8716 9004 8756
rect 9044 8716 9045 8756
rect 9003 8707 9045 8716
rect 9099 8756 9141 8765
rect 9099 8716 9100 8756
rect 9140 8716 9141 8756
rect 9099 8707 9141 8716
rect 9955 8756 10013 8757
rect 9955 8716 9964 8756
rect 10004 8716 10013 8756
rect 9955 8715 10013 8716
rect 10819 8756 10877 8757
rect 10819 8716 10828 8756
rect 10868 8716 10877 8756
rect 10819 8715 10877 8716
rect 11019 8756 11061 8765
rect 11019 8716 11020 8756
rect 11060 8716 11061 8756
rect 11019 8707 11061 8716
rect 11211 8756 11253 8765
rect 11211 8716 11212 8756
rect 11252 8716 11253 8756
rect 11211 8707 11253 8716
rect 7851 8672 7893 8681
rect 7851 8632 7852 8672
rect 7892 8632 7893 8672
rect 7851 8623 7893 8632
rect 10155 8672 10197 8681
rect 10155 8632 10156 8672
rect 10196 8632 10197 8672
rect 10155 8623 10197 8632
rect 4395 8504 4437 8513
rect 4395 8464 4396 8504
rect 4436 8464 4437 8504
rect 4395 8455 4437 8464
rect 8331 8504 8373 8513
rect 8331 8464 8332 8504
rect 8372 8464 8373 8504
rect 8331 8455 8373 8464
rect 9283 8504 9341 8505
rect 9283 8464 9292 8504
rect 9332 8464 9341 8504
rect 9283 8463 9341 8464
rect 1152 8336 11424 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 11424 8336
rect 1152 8272 11424 8296
rect 4003 8168 4061 8169
rect 4003 8128 4012 8168
rect 4052 8128 4061 8168
rect 4003 8127 4061 8128
rect 4971 8168 5013 8177
rect 4971 8128 4972 8168
rect 5012 8128 5013 8168
rect 4971 8119 5013 8128
rect 5539 8168 5597 8169
rect 5539 8128 5548 8168
rect 5588 8128 5597 8168
rect 5539 8127 5597 8128
rect 7083 8168 7125 8177
rect 7083 8128 7084 8168
rect 7124 8128 7125 8168
rect 7083 8119 7125 8128
rect 8523 8168 8565 8177
rect 8523 8128 8524 8168
rect 8564 8128 8565 8168
rect 8523 8119 8565 8128
rect 11299 8168 11357 8169
rect 11299 8128 11308 8168
rect 11348 8128 11357 8168
rect 11299 8127 11357 8128
rect 2563 7916 2621 7917
rect 2563 7876 2572 7916
rect 2612 7876 2621 7916
rect 2563 7875 2621 7876
rect 3427 7916 3485 7917
rect 3427 7876 3436 7916
rect 3476 7876 3485 7916
rect 3427 7875 3485 7876
rect 4675 7916 4733 7917
rect 4675 7876 4684 7916
rect 4724 7876 4733 7916
rect 4675 7875 4733 7876
rect 4875 7916 4917 7925
rect 4875 7876 4876 7916
rect 4916 7876 4917 7916
rect 4875 7867 4917 7876
rect 5059 7916 5117 7917
rect 5059 7876 5068 7916
rect 5108 7876 5117 7916
rect 5059 7875 5117 7876
rect 5251 7916 5309 7917
rect 5251 7876 5260 7916
rect 5300 7876 5309 7916
rect 5251 7875 5309 7876
rect 6211 7916 6269 7917
rect 6211 7876 6220 7916
rect 6260 7876 6269 7916
rect 6211 7875 6269 7876
rect 6403 7916 6461 7917
rect 6403 7876 6412 7916
rect 6452 7876 6461 7916
rect 6403 7875 6461 7876
rect 7275 7916 7317 7925
rect 7275 7876 7276 7916
rect 7316 7876 7317 7916
rect 7275 7867 7317 7876
rect 7939 7916 7997 7917
rect 7939 7876 7948 7916
rect 7988 7876 7997 7916
rect 7939 7875 7997 7876
rect 8035 7916 8093 7917
rect 8035 7876 8044 7916
rect 8084 7876 8093 7916
rect 8035 7875 8093 7876
rect 8419 7916 8477 7917
rect 8419 7876 8428 7916
rect 8468 7876 8477 7916
rect 8419 7875 8477 7876
rect 8619 7916 8661 7925
rect 8619 7876 8620 7916
rect 8660 7876 8661 7916
rect 8619 7867 8661 7876
rect 8907 7916 8949 7925
rect 8907 7876 8908 7916
rect 8948 7876 8949 7916
rect 8907 7867 8949 7876
rect 9283 7916 9341 7917
rect 9283 7876 9292 7916
rect 9332 7876 9341 7916
rect 9283 7875 9341 7876
rect 10147 7916 10205 7917
rect 10147 7876 10156 7916
rect 10196 7876 10205 7916
rect 10147 7875 10205 7876
rect 3819 7832 3861 7841
rect 3819 7792 3820 7832
rect 3860 7792 3861 7832
rect 3819 7783 3861 7792
rect 1411 7748 1469 7749
rect 1411 7708 1420 7748
rect 1460 7708 1469 7748
rect 1411 7707 1469 7708
rect 5355 7748 5397 7757
rect 5355 7708 5356 7748
rect 5396 7708 5397 7748
rect 5355 7699 5397 7708
rect 8235 7748 8277 7757
rect 8235 7708 8236 7748
rect 8276 7708 8277 7748
rect 8235 7699 8277 7708
rect 1152 7580 11424 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 11424 7580
rect 1152 7516 11424 7540
rect 1227 7412 1269 7421
rect 1227 7372 1228 7412
rect 1268 7372 1269 7412
rect 1227 7363 1269 7372
rect 3427 7412 3485 7413
rect 3427 7372 3436 7412
rect 3476 7372 3485 7412
rect 3427 7371 3485 7372
rect 4683 7412 4725 7421
rect 4683 7372 4684 7412
rect 4724 7372 4725 7412
rect 4683 7363 4725 7372
rect 6787 7412 6845 7413
rect 6787 7372 6796 7412
rect 6836 7372 6845 7412
rect 6787 7371 6845 7372
rect 9963 7412 10005 7421
rect 9963 7372 9964 7412
rect 10004 7372 10005 7412
rect 9963 7363 10005 7372
rect 1995 7328 2037 7337
rect 1995 7288 1996 7328
rect 2036 7288 2037 7328
rect 1995 7279 2037 7288
rect 9195 7328 9237 7337
rect 9195 7288 9196 7328
rect 9236 7288 9237 7328
rect 9195 7279 9237 7288
rect 1315 7244 1373 7245
rect 1315 7204 1324 7244
rect 1364 7204 1373 7244
rect 1315 7203 1373 7204
rect 1515 7244 1557 7253
rect 1515 7204 1516 7244
rect 1556 7204 1557 7244
rect 1515 7195 1557 7204
rect 1707 7244 1749 7253
rect 1707 7204 1708 7244
rect 1748 7204 1749 7244
rect 1707 7195 1749 7204
rect 1899 7244 1941 7253
rect 1899 7204 1900 7244
rect 1940 7204 1941 7244
rect 1899 7195 1941 7204
rect 2083 7244 2141 7245
rect 2083 7204 2092 7244
rect 2132 7204 2141 7244
rect 2083 7203 2141 7204
rect 2947 7244 3005 7245
rect 2947 7204 2956 7244
rect 2996 7204 3005 7244
rect 2947 7203 3005 7204
rect 3147 7244 3189 7253
rect 3147 7204 3148 7244
rect 3188 7204 3189 7244
rect 3147 7195 3189 7204
rect 3243 7244 3285 7253
rect 3243 7204 3244 7244
rect 3284 7204 3285 7244
rect 3243 7195 3285 7204
rect 3339 7244 3381 7253
rect 3339 7204 3340 7244
rect 3380 7204 3381 7244
rect 3339 7195 3381 7204
rect 3819 7244 3861 7253
rect 3819 7204 3820 7244
rect 3860 7204 3861 7244
rect 3819 7195 3861 7204
rect 4483 7244 4541 7245
rect 4483 7204 4492 7244
rect 4532 7204 4541 7244
rect 4483 7203 4541 7204
rect 4867 7244 4925 7245
rect 4867 7204 4876 7244
rect 4916 7204 4925 7244
rect 4867 7203 4925 7204
rect 4963 7244 5021 7245
rect 4963 7204 4972 7244
rect 5012 7204 5021 7244
rect 4963 7203 5021 7204
rect 5539 7244 5597 7245
rect 5539 7204 5548 7244
rect 5588 7204 5597 7244
rect 5539 7203 5597 7204
rect 7939 7244 7997 7245
rect 7939 7204 7948 7244
rect 7988 7204 7997 7244
rect 7939 7203 7997 7204
rect 8803 7244 8861 7245
rect 8803 7204 8812 7244
rect 8852 7204 8861 7244
rect 8803 7203 8861 7204
rect 10051 7244 10109 7245
rect 10051 7204 10060 7244
rect 10100 7204 10109 7244
rect 10051 7203 10109 7204
rect 10435 7244 10493 7245
rect 10435 7204 10444 7244
rect 10484 7204 10493 7244
rect 10435 7203 10493 7204
rect 10635 7244 10677 7253
rect 10635 7204 10636 7244
rect 10676 7204 10677 7244
rect 10635 7195 10677 7204
rect 11299 7244 11357 7245
rect 11299 7204 11308 7244
rect 11348 7204 11357 7244
rect 11299 7203 11357 7204
rect 1611 7160 1653 7169
rect 1611 7120 1612 7160
rect 1652 7120 1653 7160
rect 1611 7111 1653 7120
rect 5835 7076 5877 7085
rect 5835 7036 5836 7076
rect 5876 7036 5877 7076
rect 5835 7027 5877 7036
rect 2275 6992 2333 6993
rect 2275 6952 2284 6992
rect 2324 6952 2333 6992
rect 2275 6951 2333 6952
rect 6219 6992 6261 7001
rect 6219 6952 6220 6992
rect 6260 6952 6261 6992
rect 6219 6943 6261 6952
rect 1152 6824 11424 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 11424 6824
rect 1152 6760 11424 6784
rect 4483 6656 4541 6657
rect 4483 6616 4492 6656
rect 4532 6616 4541 6656
rect 4483 6615 4541 6616
rect 10923 6656 10965 6665
rect 10923 6616 10924 6656
rect 10964 6616 10965 6656
rect 10923 6607 10965 6616
rect 11115 6656 11157 6665
rect 11115 6616 11116 6656
rect 11156 6616 11157 6656
rect 11115 6607 11157 6616
rect 10155 6572 10197 6581
rect 10155 6532 10156 6572
rect 10196 6532 10197 6572
rect 10155 6523 10197 6532
rect 3627 6488 3669 6497
rect 3627 6448 3628 6488
rect 3668 6448 3669 6488
rect 3627 6439 3669 6448
rect 8323 6488 8381 6489
rect 8323 6448 8332 6488
rect 8372 6448 8381 6488
rect 8323 6447 8381 6448
rect 10723 6488 10781 6489
rect 10723 6448 10732 6488
rect 10772 6448 10781 6488
rect 10723 6447 10781 6448
rect 11299 6488 11357 6489
rect 11299 6448 11308 6488
rect 11348 6448 11357 6488
rect 11299 6447 11357 6448
rect 1227 6404 1269 6413
rect 1227 6364 1228 6404
rect 1268 6364 1269 6404
rect 1227 6355 1269 6364
rect 1603 6404 1661 6405
rect 1603 6364 1612 6404
rect 1652 6364 1661 6404
rect 1603 6363 1661 6364
rect 2467 6404 2525 6405
rect 2467 6364 2476 6404
rect 2516 6364 2525 6404
rect 2467 6363 2525 6364
rect 3811 6404 3869 6405
rect 3811 6364 3820 6404
rect 3860 6364 3869 6404
rect 3811 6363 3869 6364
rect 5059 6404 5117 6405
rect 5059 6364 5068 6404
rect 5108 6364 5117 6404
rect 5059 6363 5117 6364
rect 5923 6404 5981 6405
rect 5923 6364 5932 6404
rect 5972 6364 5981 6404
rect 5923 6363 5981 6364
rect 7363 6404 7421 6405
rect 7363 6364 7372 6404
rect 7412 6364 7421 6404
rect 7363 6363 7421 6364
rect 7563 6404 7605 6413
rect 7563 6364 7564 6404
rect 7604 6364 7605 6404
rect 7563 6355 7605 6364
rect 8035 6404 8093 6405
rect 8035 6364 8044 6404
rect 8084 6364 8093 6404
rect 8035 6363 8093 6364
rect 8131 6404 8189 6405
rect 8131 6364 8140 6404
rect 8180 6364 8189 6404
rect 8131 6363 8189 6364
rect 9475 6404 9533 6405
rect 9475 6364 9484 6404
rect 9524 6364 9533 6404
rect 9475 6363 9533 6364
rect 4683 6320 4725 6329
rect 4683 6280 4684 6320
rect 4724 6280 4725 6320
rect 4683 6271 4725 6280
rect 7467 6320 7509 6329
rect 7467 6280 7468 6320
rect 7508 6280 7509 6320
rect 7467 6271 7509 6280
rect 7075 6236 7133 6237
rect 7075 6196 7084 6236
rect 7124 6196 7133 6236
rect 7075 6195 7133 6196
rect 1152 6068 11424 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 11424 6068
rect 1152 6004 11424 6028
rect 1419 5900 1461 5909
rect 1419 5860 1420 5900
rect 1460 5860 1461 5900
rect 1419 5851 1461 5860
rect 1803 5900 1845 5909
rect 1803 5860 1804 5900
rect 1844 5860 1845 5900
rect 1803 5851 1845 5860
rect 3819 5900 3861 5909
rect 3819 5860 3820 5900
rect 3860 5860 3861 5900
rect 3819 5851 3861 5860
rect 11203 5900 11261 5901
rect 11203 5860 11212 5900
rect 11252 5860 11261 5900
rect 11203 5859 11261 5860
rect 8811 5816 8853 5825
rect 8811 5776 8812 5816
rect 8852 5776 8853 5816
rect 8811 5767 8853 5776
rect 1995 5732 2037 5741
rect 1995 5692 1996 5732
rect 2036 5692 2037 5732
rect 1995 5683 2037 5692
rect 2083 5732 2141 5733
rect 2083 5692 2092 5732
rect 2132 5692 2141 5732
rect 2083 5691 2141 5692
rect 2475 5732 2517 5741
rect 2475 5692 2476 5732
rect 2516 5692 2517 5732
rect 2475 5683 2517 5692
rect 2571 5732 2613 5741
rect 2571 5692 2572 5732
rect 2612 5692 2613 5732
rect 2571 5683 2613 5692
rect 2659 5732 2717 5733
rect 2659 5692 2668 5732
rect 2708 5692 2717 5732
rect 2659 5691 2717 5692
rect 2859 5732 2901 5741
rect 2859 5692 2860 5732
rect 2900 5692 2901 5732
rect 2859 5683 2901 5692
rect 3043 5732 3101 5733
rect 3043 5692 3052 5732
rect 3092 5692 3101 5732
rect 3043 5691 3101 5692
rect 3435 5732 3477 5741
rect 3435 5692 3436 5732
rect 3476 5692 3477 5732
rect 3435 5683 3477 5692
rect 3523 5732 3581 5733
rect 3523 5692 3532 5732
rect 3572 5692 3581 5732
rect 3523 5691 3581 5692
rect 4875 5732 4917 5741
rect 4875 5692 4876 5732
rect 4916 5692 4917 5732
rect 4875 5683 4917 5692
rect 5923 5732 5981 5733
rect 5923 5692 5932 5732
rect 5972 5692 5981 5732
rect 5923 5691 5981 5692
rect 6211 5732 6269 5733
rect 6211 5692 6220 5732
rect 6260 5692 6269 5732
rect 6211 5691 6269 5692
rect 7075 5732 7133 5733
rect 7075 5692 7084 5732
rect 7124 5692 7133 5732
rect 7075 5691 7133 5692
rect 7939 5732 7997 5733
rect 7939 5692 7948 5732
rect 7988 5692 7997 5732
rect 7939 5691 7997 5692
rect 8131 5732 8189 5733
rect 8131 5692 8140 5732
rect 8180 5692 8189 5732
rect 8131 5691 8189 5692
rect 8235 5732 8277 5741
rect 8235 5692 8236 5732
rect 8276 5692 8277 5732
rect 8235 5683 8277 5692
rect 8427 5732 8469 5741
rect 8427 5692 8428 5732
rect 8468 5692 8469 5732
rect 8427 5683 8469 5692
rect 8619 5732 8661 5741
rect 8619 5692 8620 5732
rect 8660 5692 8661 5732
rect 8619 5683 8661 5692
rect 9187 5732 9245 5733
rect 9187 5692 9196 5732
rect 9236 5692 9245 5732
rect 9187 5691 9245 5692
rect 10051 5732 10109 5733
rect 10051 5692 10060 5732
rect 10100 5692 10109 5732
rect 10051 5691 10109 5692
rect 1219 5648 1277 5649
rect 1219 5608 1228 5648
rect 1268 5608 1277 5648
rect 1219 5607 1277 5608
rect 1603 5648 1661 5649
rect 1603 5608 1612 5648
rect 1652 5608 1661 5648
rect 1603 5607 1661 5608
rect 2955 5648 2997 5657
rect 2955 5608 2956 5648
rect 2996 5608 2997 5648
rect 2955 5599 2997 5608
rect 4683 5480 4725 5489
rect 4683 5440 4684 5480
rect 4724 5440 4725 5480
rect 4683 5431 4725 5440
rect 5251 5480 5309 5481
rect 5251 5440 5260 5480
rect 5300 5440 5309 5480
rect 5251 5439 5309 5440
rect 6123 5480 6165 5489
rect 6123 5440 6124 5480
rect 6164 5440 6165 5480
rect 6123 5431 6165 5440
rect 6403 5480 6461 5481
rect 6403 5440 6412 5480
rect 6452 5440 6461 5480
rect 6403 5439 6461 5440
rect 7267 5480 7325 5481
rect 7267 5440 7276 5480
rect 7316 5440 7325 5480
rect 7267 5439 7325 5440
rect 8427 5480 8469 5489
rect 8427 5440 8428 5480
rect 8468 5440 8469 5480
rect 8427 5431 8469 5440
rect 1152 5312 11424 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 11424 5312
rect 1152 5248 11424 5272
rect 8323 5060 8381 5061
rect 8323 5020 8332 5060
rect 8372 5020 8381 5060
rect 8323 5019 8381 5020
rect 11115 5060 11157 5069
rect 11115 5020 11116 5060
rect 11156 5020 11157 5060
rect 11115 5011 11157 5020
rect 11299 4976 11357 4977
rect 11299 4936 11308 4976
rect 11348 4936 11357 4976
rect 11299 4935 11357 4936
rect 2763 4892 2805 4901
rect 2763 4852 2764 4892
rect 2804 4852 2805 4892
rect 2763 4843 2805 4852
rect 2955 4892 2997 4901
rect 2955 4852 2956 4892
rect 2996 4852 2997 4892
rect 2955 4843 2997 4852
rect 3147 4892 3189 4901
rect 3147 4852 3148 4892
rect 3188 4852 3189 4892
rect 3147 4843 3189 4852
rect 3243 4892 3285 4901
rect 3243 4852 3244 4892
rect 3284 4852 3285 4892
rect 3243 4843 3285 4852
rect 3339 4892 3381 4901
rect 3339 4852 3340 4892
rect 3380 4852 3381 4892
rect 3339 4843 3381 4852
rect 3435 4892 3477 4901
rect 3435 4852 3436 4892
rect 3476 4852 3477 4892
rect 3435 4843 3477 4852
rect 4291 4892 4349 4893
rect 4291 4852 4300 4892
rect 4340 4852 4349 4892
rect 4291 4851 4349 4852
rect 4771 4892 4829 4893
rect 4771 4852 4780 4892
rect 4820 4852 4829 4892
rect 4771 4851 4829 4852
rect 4867 4892 4925 4893
rect 4867 4852 4876 4892
rect 4916 4852 4925 4892
rect 4867 4851 4925 4852
rect 5251 4892 5309 4893
rect 5251 4852 5260 4892
rect 5300 4852 5309 4892
rect 5251 4851 5309 4852
rect 6115 4892 6173 4893
rect 6115 4852 6124 4892
rect 6164 4852 6173 4892
rect 6115 4851 6173 4852
rect 6403 4892 6461 4893
rect 6403 4852 6412 4892
rect 6452 4852 6461 4892
rect 6403 4851 6461 4852
rect 6691 4892 6749 4893
rect 6691 4852 6700 4892
rect 6740 4852 6749 4892
rect 6691 4851 6749 4852
rect 7843 4892 7901 4893
rect 7843 4852 7852 4892
rect 7892 4852 7901 4892
rect 7843 4851 7901 4852
rect 8995 4892 9053 4893
rect 8995 4852 9004 4892
rect 9044 4852 9053 4892
rect 8995 4851 9053 4852
rect 5931 4808 5973 4817
rect 5931 4768 5932 4808
rect 5972 4768 5973 4808
rect 5931 4759 5973 4768
rect 6883 4808 6941 4809
rect 6883 4768 6892 4808
rect 6932 4768 6941 4808
rect 6883 4767 6941 4768
rect 2859 4724 2901 4733
rect 2859 4684 2860 4724
rect 2900 4684 2901 4724
rect 2859 4675 2901 4684
rect 3619 4724 3677 4725
rect 3619 4684 3628 4724
rect 3668 4684 3677 4724
rect 3619 4683 3677 4684
rect 5067 4724 5109 4733
rect 5067 4684 5068 4724
rect 5108 4684 5109 4724
rect 5067 4675 5109 4684
rect 6219 4724 6261 4733
rect 6219 4684 6220 4724
rect 6260 4684 6261 4724
rect 6219 4675 6261 4684
rect 7171 4724 7229 4725
rect 7171 4684 7180 4724
rect 7220 4684 7229 4724
rect 7171 4683 7229 4684
rect 1152 4556 11424 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 11424 4556
rect 1152 4492 11424 4516
rect 5059 4388 5117 4389
rect 5059 4348 5068 4388
rect 5108 4348 5117 4388
rect 5059 4347 5117 4348
rect 6595 4388 6653 4389
rect 6595 4348 6604 4388
rect 6644 4348 6653 4388
rect 6595 4347 6653 4348
rect 9475 4388 9533 4389
rect 9475 4348 9484 4388
rect 9524 4348 9533 4388
rect 9475 4347 9533 4348
rect 2667 4304 2709 4313
rect 2667 4264 2668 4304
rect 2708 4264 2709 4304
rect 2667 4255 2709 4264
rect 5347 4304 5405 4305
rect 5347 4264 5356 4304
rect 5396 4264 5405 4304
rect 5347 4263 5405 4264
rect 6315 4304 6357 4313
rect 6315 4264 6316 4304
rect 6356 4264 6357 4304
rect 6315 4255 6357 4264
rect 3043 4220 3101 4221
rect 3043 4180 3052 4220
rect 3092 4180 3101 4220
rect 3043 4179 3101 4180
rect 3907 4220 3965 4221
rect 3907 4180 3916 4220
rect 3956 4180 3965 4220
rect 3907 4179 3965 4180
rect 5443 4220 5501 4221
rect 5443 4180 5452 4220
rect 5492 4180 5501 4220
rect 5443 4179 5501 4180
rect 5827 4220 5885 4221
rect 5827 4180 5836 4220
rect 5876 4180 5885 4220
rect 5827 4179 5885 4180
rect 6219 4220 6261 4229
rect 6219 4180 6220 4220
rect 6260 4180 6261 4220
rect 6219 4171 6261 4180
rect 6403 4220 6461 4221
rect 6403 4180 6412 4220
rect 6452 4180 6461 4220
rect 6403 4179 6461 4180
rect 6699 4220 6741 4229
rect 6699 4180 6700 4220
rect 6740 4180 6741 4220
rect 6699 4171 6741 4180
rect 6795 4220 6837 4229
rect 6795 4180 6796 4220
rect 6836 4180 6837 4220
rect 6795 4171 6837 4180
rect 6891 4220 6933 4229
rect 6891 4180 6892 4220
rect 6932 4180 6933 4220
rect 6891 4171 6933 4180
rect 7083 4220 7125 4229
rect 7083 4180 7084 4220
rect 7124 4180 7125 4220
rect 7083 4171 7125 4180
rect 7459 4220 7517 4221
rect 7459 4180 7468 4220
rect 7508 4180 7517 4220
rect 7459 4179 7517 4180
rect 8323 4220 8381 4221
rect 8323 4180 8332 4220
rect 8372 4180 8381 4220
rect 8323 4179 8381 4180
rect 1152 3800 11424 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 11424 3800
rect 1152 3736 11424 3760
rect 3147 3632 3189 3641
rect 3147 3592 3148 3632
rect 3188 3592 3189 3632
rect 3147 3583 3189 3592
rect 5163 3632 5205 3641
rect 5163 3592 5164 3632
rect 5204 3592 5205 3632
rect 5163 3583 5205 3592
rect 7843 3632 7901 3633
rect 7843 3592 7852 3632
rect 7892 3592 7901 3632
rect 7843 3591 7901 3592
rect 8035 3632 8093 3633
rect 8035 3592 8044 3632
rect 8084 3592 8093 3632
rect 8035 3591 8093 3592
rect 8907 3548 8949 3557
rect 8907 3508 8908 3548
rect 8948 3508 8949 3548
rect 8907 3499 8949 3508
rect 9091 3464 9149 3465
rect 9091 3424 9100 3464
rect 9140 3424 9149 3464
rect 9091 3423 9149 3424
rect 3235 3380 3293 3381
rect 3235 3340 3244 3380
rect 3284 3340 3293 3380
rect 3235 3339 3293 3340
rect 5059 3380 5117 3381
rect 5059 3340 5068 3380
rect 5108 3340 5117 3380
rect 5059 3339 5117 3340
rect 5259 3380 5301 3389
rect 5259 3340 5260 3380
rect 5300 3340 5301 3380
rect 5259 3331 5301 3340
rect 5451 3380 5493 3389
rect 5451 3340 5452 3380
rect 5492 3340 5493 3380
rect 5451 3331 5493 3340
rect 5827 3380 5885 3381
rect 5827 3340 5836 3380
rect 5876 3340 5885 3380
rect 5827 3339 5885 3340
rect 6691 3380 6749 3381
rect 6691 3340 6700 3380
rect 6740 3340 6749 3380
rect 6691 3339 6749 3340
rect 8707 3380 8765 3381
rect 8707 3340 8716 3380
rect 8756 3340 8765 3380
rect 8707 3339 8765 3340
rect 1152 3044 11424 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 11424 3044
rect 1152 2980 11424 3004
<< via1 >>
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 2860 12496 2900 12536
rect 7468 12496 7508 12536
rect 3244 12412 3284 12452
rect 3628 12412 3668 12452
rect 4684 12412 4724 12452
rect 4876 12412 4916 12452
rect 5068 12412 5108 12452
rect 5356 12412 5396 12452
rect 6028 12412 6068 12452
rect 6316 12412 6356 12452
rect 8716 12412 8756 12452
rect 4972 12328 5012 12368
rect 3052 12244 3092 12284
rect 3724 12244 3764 12284
rect 4012 12244 4052 12284
rect 6412 12244 6452 12284
rect 7276 12244 7316 12284
rect 9388 12244 9428 12284
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 1900 11908 1940 11948
rect 5932 11908 5972 11948
rect 8524 11908 8564 11948
rect 3532 11824 3572 11864
rect 1228 11740 1268 11780
rect 1420 11740 1460 11780
rect 2188 11740 2228 11780
rect 2860 11740 2900 11780
rect 3148 11740 3188 11780
rect 3340 11740 3380 11780
rect 3916 11740 3956 11780
rect 4780 11740 4820 11780
rect 6124 11740 6164 11780
rect 6508 11740 6548 11780
rect 7372 11740 7412 11780
rect 9388 11740 9428 11780
rect 9580 11740 9620 11780
rect 9772 11740 9812 11780
rect 10636 11740 10676 11780
rect 1708 11656 1748 11696
rect 2956 11656 2996 11696
rect 9676 11572 9716 11612
rect 2092 11488 2132 11528
rect 3340 11488 3380 11528
rect 8716 11488 8756 11528
rect 9964 11488 10004 11528
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 11116 11152 11156 11192
rect 5836 10984 5876 11024
rect 1996 10900 2036 10940
rect 2860 10900 2900 10940
rect 4396 10900 4436 10940
rect 5452 10900 5492 10940
rect 5548 10900 5588 10940
rect 6412 10900 6452 10940
rect 7564 10900 7604 10940
rect 7756 10900 7796 10940
rect 8236 10900 8276 10940
rect 8524 10900 8564 10940
rect 9100 10900 9140 10940
rect 9964 10900 10004 10940
rect 1612 10816 1652 10856
rect 8716 10816 8756 10856
rect 4012 10732 4052 10772
rect 5068 10732 5108 10772
rect 6892 10732 6932 10772
rect 7660 10732 7700 10772
rect 8044 10732 8084 10772
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 1324 10396 1364 10436
rect 3436 10396 3476 10436
rect 4876 10396 4916 10436
rect 5068 10396 5108 10436
rect 5836 10396 5876 10436
rect 8812 10396 8852 10436
rect 9964 10312 10004 10352
rect 1516 10228 1556 10268
rect 1612 10228 1652 10268
rect 2764 10228 2804 10268
rect 2956 10228 2996 10268
rect 3916 10228 3956 10268
rect 4204 10228 4244 10268
rect 5164 10228 5204 10268
rect 5260 10228 5300 10268
rect 5356 10228 5396 10268
rect 5548 10228 5588 10268
rect 5644 10228 5684 10268
rect 5740 10228 5780 10268
rect 6124 10228 6164 10268
rect 6988 10228 7028 10268
rect 7180 10228 7220 10268
rect 7660 10228 7700 10268
rect 7756 10228 7796 10268
rect 8140 10228 8180 10268
rect 9196 10228 9236 10268
rect 10252 10228 10292 10268
rect 10444 10228 10484 10268
rect 11308 10228 11348 10268
rect 7084 10144 7124 10184
rect 7948 10144 7988 10184
rect 2092 10060 2132 10100
rect 9388 10060 9428 10100
rect 10636 10060 10676 10100
rect 6028 9976 6068 10016
rect 9772 9976 9812 10016
rect 10348 9976 10388 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 4012 9640 4052 9680
rect 4396 9640 4436 9680
rect 11020 9640 11060 9680
rect 1228 9472 1268 9512
rect 1996 9388 2036 9428
rect 2860 9388 2900 9428
rect 4300 9388 4340 9428
rect 4492 9388 4532 9428
rect 4684 9388 4724 9428
rect 5068 9388 5108 9428
rect 6220 9388 6260 9428
rect 6412 9388 6452 9428
rect 6604 9388 6644 9428
rect 6796 9388 6836 9428
rect 7468 9388 7508 9428
rect 7852 9388 7892 9428
rect 8140 9388 8180 9428
rect 8236 9388 8276 9428
rect 8332 9388 8372 9428
rect 8428 9388 8468 9428
rect 8620 9388 8660 9428
rect 9004 9388 9044 9428
rect 9868 9388 9908 9428
rect 1612 9304 1652 9344
rect 6508 9304 6548 9344
rect 1420 9220 1460 9260
rect 5164 9220 5204 9260
rect 5548 9220 5588 9260
rect 7948 9220 7988 9260
rect 11020 9220 11060 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 1996 8884 2036 8924
rect 5260 8884 5300 8924
rect 2860 8800 2900 8840
rect 3244 8800 3284 8840
rect 3628 8800 3668 8840
rect 5452 8800 5492 8840
rect 8620 8800 8660 8840
rect 11116 8800 11156 8840
rect 1708 8716 1748 8756
rect 1804 8716 1844 8756
rect 2188 8716 2228 8756
rect 2284 8716 2324 8756
rect 2764 8716 2804 8756
rect 2956 8716 2996 8756
rect 3148 8716 3188 8756
rect 3340 8716 3380 8756
rect 3820 8716 3860 8756
rect 4108 8716 4148 8756
rect 4300 8716 4340 8756
rect 4588 8716 4628 8756
rect 5836 8716 5876 8756
rect 6700 8716 6740 8756
rect 8236 8716 8276 8756
rect 8524 8716 8564 8756
rect 8812 8716 8852 8756
rect 8908 8716 8948 8756
rect 9004 8716 9044 8756
rect 9100 8716 9140 8756
rect 9964 8716 10004 8756
rect 10828 8716 10868 8756
rect 11020 8716 11060 8756
rect 11212 8716 11252 8756
rect 7852 8632 7892 8672
rect 10156 8632 10196 8672
rect 4396 8464 4436 8504
rect 8332 8464 8372 8504
rect 9292 8464 9332 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4012 8128 4052 8168
rect 4972 8128 5012 8168
rect 5548 8128 5588 8168
rect 7084 8128 7124 8168
rect 8524 8128 8564 8168
rect 11308 8128 11348 8168
rect 2572 7876 2612 7916
rect 3436 7876 3476 7916
rect 4684 7876 4724 7916
rect 4876 7876 4916 7916
rect 5068 7876 5108 7916
rect 5260 7876 5300 7916
rect 6220 7876 6260 7916
rect 6412 7876 6452 7916
rect 7276 7876 7316 7916
rect 7948 7876 7988 7916
rect 8044 7876 8084 7916
rect 8428 7876 8468 7916
rect 8620 7876 8660 7916
rect 8908 7876 8948 7916
rect 9292 7876 9332 7916
rect 10156 7876 10196 7916
rect 3820 7792 3860 7832
rect 1420 7708 1460 7748
rect 5356 7708 5396 7748
rect 8236 7708 8276 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 1228 7372 1268 7412
rect 3436 7372 3476 7412
rect 4684 7372 4724 7412
rect 6796 7372 6836 7412
rect 9964 7372 10004 7412
rect 1996 7288 2036 7328
rect 9196 7288 9236 7328
rect 1324 7204 1364 7244
rect 1516 7204 1556 7244
rect 1708 7204 1748 7244
rect 1900 7204 1940 7244
rect 2092 7204 2132 7244
rect 2956 7204 2996 7244
rect 3148 7204 3188 7244
rect 3244 7204 3284 7244
rect 3340 7204 3380 7244
rect 3820 7204 3860 7244
rect 4492 7204 4532 7244
rect 4876 7204 4916 7244
rect 4972 7204 5012 7244
rect 5548 7204 5588 7244
rect 7948 7204 7988 7244
rect 8812 7204 8852 7244
rect 10060 7204 10100 7244
rect 10444 7204 10484 7244
rect 10636 7204 10676 7244
rect 11308 7204 11348 7244
rect 1612 7120 1652 7160
rect 5836 7036 5876 7076
rect 2284 6952 2324 6992
rect 6220 6952 6260 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4492 6616 4532 6656
rect 10924 6616 10964 6656
rect 11116 6616 11156 6656
rect 10156 6532 10196 6572
rect 3628 6448 3668 6488
rect 8332 6448 8372 6488
rect 10732 6448 10772 6488
rect 11308 6448 11348 6488
rect 1228 6364 1268 6404
rect 1612 6364 1652 6404
rect 2476 6364 2516 6404
rect 3820 6364 3860 6404
rect 5068 6364 5108 6404
rect 5932 6364 5972 6404
rect 7372 6364 7412 6404
rect 7564 6364 7604 6404
rect 8044 6364 8084 6404
rect 8140 6364 8180 6404
rect 9484 6364 9524 6404
rect 4684 6280 4724 6320
rect 7468 6280 7508 6320
rect 7084 6196 7124 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 1420 5860 1460 5900
rect 1804 5860 1844 5900
rect 3820 5860 3860 5900
rect 11212 5860 11252 5900
rect 8812 5776 8852 5816
rect 1996 5692 2036 5732
rect 2092 5692 2132 5732
rect 2476 5692 2516 5732
rect 2572 5692 2612 5732
rect 2668 5692 2708 5732
rect 2860 5692 2900 5732
rect 3052 5692 3092 5732
rect 3436 5692 3476 5732
rect 3532 5692 3572 5732
rect 4876 5692 4916 5732
rect 5932 5692 5972 5732
rect 6220 5692 6260 5732
rect 7084 5692 7124 5732
rect 7948 5692 7988 5732
rect 8140 5692 8180 5732
rect 8236 5692 8276 5732
rect 8428 5692 8468 5732
rect 8620 5692 8660 5732
rect 9196 5692 9236 5732
rect 10060 5692 10100 5732
rect 1228 5608 1268 5648
rect 1612 5608 1652 5648
rect 2956 5608 2996 5648
rect 4684 5440 4724 5480
rect 5260 5440 5300 5480
rect 6124 5440 6164 5480
rect 6412 5440 6452 5480
rect 7276 5440 7316 5480
rect 8428 5440 8468 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 8332 5020 8372 5060
rect 11116 5020 11156 5060
rect 11308 4936 11348 4976
rect 2764 4852 2804 4892
rect 2956 4852 2996 4892
rect 3148 4852 3188 4892
rect 3244 4852 3284 4892
rect 3340 4852 3380 4892
rect 3436 4852 3476 4892
rect 4300 4852 4340 4892
rect 4780 4852 4820 4892
rect 4876 4852 4916 4892
rect 5260 4852 5300 4892
rect 6124 4852 6164 4892
rect 6412 4852 6452 4892
rect 6700 4852 6740 4892
rect 7852 4852 7892 4892
rect 9004 4852 9044 4892
rect 5932 4768 5972 4808
rect 6892 4768 6932 4808
rect 2860 4684 2900 4724
rect 3628 4684 3668 4724
rect 5068 4684 5108 4724
rect 6220 4684 6260 4724
rect 7180 4684 7220 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 5068 4348 5108 4388
rect 6604 4348 6644 4388
rect 9484 4348 9524 4388
rect 2668 4264 2708 4304
rect 5356 4264 5396 4304
rect 6316 4264 6356 4304
rect 3052 4180 3092 4220
rect 3916 4180 3956 4220
rect 5452 4180 5492 4220
rect 5836 4180 5876 4220
rect 6220 4180 6260 4220
rect 6412 4180 6452 4220
rect 6700 4180 6740 4220
rect 6796 4180 6836 4220
rect 6892 4180 6932 4220
rect 7084 4180 7124 4220
rect 7468 4180 7508 4220
rect 8332 4180 8372 4220
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 3148 3592 3188 3632
rect 5164 3592 5204 3632
rect 7852 3592 7892 3632
rect 8044 3592 8084 3632
rect 8908 3508 8948 3548
rect 9100 3424 9140 3464
rect 3244 3340 3284 3380
rect 5068 3340 5108 3380
rect 5260 3340 5300 3380
rect 5452 3340 5492 3380
rect 5836 3340 5876 3380
rect 6700 3340 6740 3380
rect 8716 3340 8756 3380
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
<< metal2 >>
rect 4088 16248 4168 16328
rect 7160 16248 7240 16328
rect 4108 13889 4148 16248
rect 2859 13880 2901 13889
rect 2859 13840 2860 13880
rect 2900 13840 2901 13880
rect 2859 13831 2901 13840
rect 4107 13880 4149 13889
rect 4107 13840 4108 13880
rect 4148 13840 4149 13880
rect 4107 13831 4149 13840
rect 2860 12536 2900 13831
rect 3688 12872 4056 12881
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 3688 12823 4056 12832
rect 3147 12620 3189 12629
rect 3147 12580 3148 12620
rect 3188 12580 3189 12620
rect 3147 12571 3189 12580
rect 5067 12620 5109 12629
rect 5067 12580 5068 12620
rect 5108 12580 5109 12620
rect 5067 12571 5109 12580
rect 5931 12620 5973 12629
rect 5931 12580 5932 12620
rect 5972 12580 5973 12620
rect 5931 12571 5973 12580
rect 2860 12487 2900 12496
rect 3052 12284 3092 12293
rect 3052 11957 3092 12244
rect 1899 11948 1941 11957
rect 1899 11908 1900 11948
rect 1940 11908 1941 11948
rect 1899 11899 1941 11908
rect 3051 11948 3093 11957
rect 3051 11908 3052 11948
rect 3092 11908 3093 11948
rect 3051 11899 3093 11908
rect 1900 11814 1940 11899
rect 1228 11780 1268 11789
rect 1228 11369 1268 11740
rect 1420 11780 1460 11789
rect 1420 11369 1460 11740
rect 2188 11780 2228 11789
rect 2379 11780 2421 11789
rect 2228 11740 2380 11780
rect 2420 11740 2421 11780
rect 2188 11731 2228 11740
rect 2379 11731 2421 11740
rect 2859 11780 2901 11789
rect 2859 11740 2860 11780
rect 2900 11740 2901 11780
rect 2859 11731 2901 11740
rect 3148 11780 3188 12571
rect 3339 12536 3381 12545
rect 3339 12496 3340 12536
rect 3380 12496 3381 12536
rect 3339 12487 3381 12496
rect 3627 12536 3669 12545
rect 3627 12496 3628 12536
rect 3668 12496 3669 12536
rect 3627 12487 3669 12496
rect 4587 12536 4629 12545
rect 4587 12496 4588 12536
rect 4628 12496 4629 12536
rect 4587 12487 4629 12496
rect 4875 12536 4917 12545
rect 4875 12496 4876 12536
rect 4916 12496 4917 12536
rect 4875 12487 4917 12496
rect 3243 12452 3285 12461
rect 3243 12412 3244 12452
rect 3284 12412 3285 12452
rect 3243 12403 3285 12412
rect 3244 12318 3284 12403
rect 3148 11731 3188 11740
rect 3340 11780 3380 12487
rect 3628 12452 3668 12487
rect 3628 12401 3668 12412
rect 4395 12368 4437 12377
rect 4395 12328 4396 12368
rect 4436 12328 4437 12368
rect 4395 12319 4437 12328
rect 3724 12284 3764 12293
rect 3819 12284 3861 12293
rect 3764 12244 3820 12284
rect 3860 12244 3861 12284
rect 3724 12235 3764 12244
rect 3819 12235 3861 12244
rect 4012 12284 4052 12293
rect 4012 11873 4052 12244
rect 4299 11948 4341 11957
rect 4299 11908 4300 11948
rect 4340 11908 4341 11948
rect 4299 11899 4341 11908
rect 3531 11864 3573 11873
rect 3531 11824 3532 11864
rect 3572 11824 3573 11864
rect 3531 11815 3573 11824
rect 4011 11864 4053 11873
rect 4011 11824 4012 11864
rect 4052 11824 4053 11864
rect 4011 11815 4053 11824
rect 3340 11731 3380 11740
rect 3435 11780 3477 11789
rect 3435 11740 3436 11780
rect 3476 11740 3477 11780
rect 3435 11731 3477 11740
rect 1708 11696 1748 11705
rect 1708 11537 1748 11656
rect 1707 11528 1749 11537
rect 1707 11488 1708 11528
rect 1748 11488 1749 11528
rect 1707 11479 1749 11488
rect 2092 11528 2132 11537
rect 1227 11360 1269 11369
rect 1227 11320 1228 11360
rect 1268 11320 1269 11360
rect 1227 11311 1269 11320
rect 1419 11360 1461 11369
rect 2092 11360 2132 11488
rect 1419 11320 1420 11360
rect 1460 11320 1461 11360
rect 1419 11311 1461 11320
rect 1996 11320 2132 11360
rect 1996 10940 2036 11320
rect 1996 10891 2036 10900
rect 1612 10856 1652 10865
rect 1324 10816 1612 10856
rect 1324 10436 1364 10816
rect 1612 10807 1652 10816
rect 1324 10387 1364 10396
rect 1516 10268 1556 10277
rect 1228 9512 1268 9521
rect 1228 9185 1268 9472
rect 1420 9260 1460 9269
rect 1227 9176 1269 9185
rect 1227 9136 1228 9176
rect 1268 9136 1269 9176
rect 1227 9127 1269 9136
rect 1420 8765 1460 9220
rect 1516 8849 1556 10228
rect 1612 10268 1652 10277
rect 1612 10100 1652 10228
rect 2092 10100 2132 10109
rect 1612 10060 2092 10100
rect 2132 10060 2324 10100
rect 2092 10051 2132 10060
rect 1996 9428 2036 9437
rect 2036 9388 2132 9428
rect 1996 9379 2036 9388
rect 1612 9344 1652 9353
rect 1652 9304 1844 9344
rect 1612 9295 1652 9304
rect 1804 8924 1844 9304
rect 1996 8924 2036 8933
rect 1804 8884 1996 8924
rect 1996 8875 2036 8884
rect 1515 8840 1557 8849
rect 1515 8800 1516 8840
rect 1556 8800 1557 8840
rect 1515 8791 1557 8800
rect 1419 8756 1461 8765
rect 1419 8716 1420 8756
rect 1460 8716 1461 8756
rect 1419 8707 1461 8716
rect 1708 8756 1748 8767
rect 1708 8681 1748 8716
rect 1804 8756 1844 8765
rect 2092 8756 2132 9388
rect 2187 8840 2229 8849
rect 2187 8800 2188 8840
rect 2228 8800 2229 8840
rect 2187 8791 2229 8800
rect 1844 8716 2132 8756
rect 2188 8756 2228 8791
rect 1804 8707 1844 8716
rect 2188 8705 2228 8716
rect 2284 8756 2324 10060
rect 2284 8707 2324 8716
rect 2380 8681 2420 11731
rect 2860 11646 2900 11731
rect 2955 11696 2997 11705
rect 2955 11656 2956 11696
rect 2996 11656 2997 11696
rect 2955 11647 2997 11656
rect 2956 11562 2996 11647
rect 3340 11528 3380 11537
rect 2955 11360 2997 11369
rect 2955 11320 2956 11360
rect 2996 11320 3092 11360
rect 2955 11311 2997 11320
rect 2860 10940 2900 10949
rect 2764 10268 2804 10277
rect 2764 10109 2804 10228
rect 2860 10268 2900 10900
rect 2956 10268 2996 10277
rect 2860 10228 2956 10268
rect 2763 10100 2805 10109
rect 2763 10060 2764 10100
rect 2804 10060 2805 10100
rect 2763 10051 2805 10060
rect 2860 9428 2900 10228
rect 2956 10219 2996 10228
rect 3052 9521 3092 11320
rect 3340 10193 3380 11488
rect 3436 10436 3476 11731
rect 3532 11730 3572 11815
rect 3916 11780 3956 11791
rect 3916 11705 3956 11740
rect 3915 11696 3957 11705
rect 3915 11656 3916 11696
rect 3956 11656 3957 11696
rect 3915 11647 3957 11656
rect 3688 11360 4056 11369
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 3688 11311 4056 11320
rect 4012 10772 4052 10781
rect 4052 10732 4244 10772
rect 4012 10723 4052 10732
rect 3436 10387 3476 10396
rect 3916 10268 3956 10277
rect 4204 10268 4244 10732
rect 3956 10228 4148 10268
rect 3916 10219 3956 10228
rect 3339 10184 3381 10193
rect 3339 10144 3340 10184
rect 3380 10144 3381 10184
rect 3339 10135 3381 10144
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 4011 9680 4053 9689
rect 4011 9640 4012 9680
rect 4052 9640 4053 9680
rect 4011 9631 4053 9640
rect 4012 9546 4052 9631
rect 3051 9512 3093 9521
rect 3051 9472 3052 9512
rect 3092 9472 3093 9512
rect 3051 9463 3093 9472
rect 2668 9388 2860 9428
rect 1323 8672 1365 8681
rect 1323 8632 1324 8672
rect 1364 8632 1365 8672
rect 1323 8623 1365 8632
rect 1707 8672 1749 8681
rect 1707 8632 1708 8672
rect 1748 8632 1749 8672
rect 1707 8623 1749 8632
rect 2379 8672 2421 8681
rect 2379 8632 2380 8672
rect 2420 8632 2421 8672
rect 2379 8623 2421 8632
rect 1227 7580 1269 7589
rect 1227 7540 1228 7580
rect 1268 7540 1269 7580
rect 1227 7531 1269 7540
rect 1228 7412 1268 7531
rect 1228 7363 1268 7372
rect 1324 7244 1364 8623
rect 2572 7916 2612 7925
rect 2668 7916 2708 9388
rect 2860 9379 2900 9388
rect 2859 8840 2901 8849
rect 2859 8800 2860 8840
rect 2900 8800 2901 8840
rect 2859 8791 2901 8800
rect 2763 8756 2805 8765
rect 2763 8716 2764 8756
rect 2804 8716 2805 8756
rect 2763 8707 2805 8716
rect 2764 8622 2804 8707
rect 2860 8706 2900 8791
rect 2956 8756 2996 8765
rect 3052 8756 3092 9463
rect 3147 9428 3189 9437
rect 3147 9388 3148 9428
rect 3188 9388 3189 9428
rect 3147 9379 3189 9388
rect 2996 8716 3092 8756
rect 3148 8756 3188 9379
rect 4108 8924 4148 10228
rect 4204 10219 4244 10228
rect 4300 9428 4340 11899
rect 4396 10940 4436 12319
rect 4396 10891 4436 10900
rect 4588 10688 4628 12487
rect 4684 12452 4724 12461
rect 4684 11360 4724 12412
rect 4876 12452 4916 12487
rect 4876 12401 4916 12412
rect 4972 12377 5012 12462
rect 5068 12452 5108 12571
rect 5068 12403 5108 12412
rect 5355 12452 5397 12461
rect 5355 12412 5356 12452
rect 5396 12412 5397 12452
rect 5355 12403 5397 12412
rect 5932 12452 5972 12571
rect 7180 12536 7220 16248
rect 7468 12536 7508 12545
rect 7180 12496 7468 12536
rect 7468 12487 7508 12496
rect 6028 12452 6068 12480
rect 5932 12412 6028 12452
rect 4971 12368 5013 12377
rect 4971 12328 4972 12368
rect 5012 12328 5013 12368
rect 4971 12319 5013 12328
rect 5356 12318 5396 12403
rect 5451 12284 5493 12293
rect 5451 12244 5452 12284
rect 5492 12244 5493 12284
rect 5451 12235 5493 12244
rect 4928 12116 5296 12125
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 4928 12067 5296 12076
rect 4779 11780 4821 11789
rect 4779 11740 4780 11780
rect 4820 11740 4821 11780
rect 4779 11731 4821 11740
rect 4780 11646 4820 11731
rect 4684 11320 4820 11360
rect 4588 10648 4724 10688
rect 4684 10436 4724 10648
rect 4780 10613 4820 11320
rect 5452 10940 5492 12235
rect 5932 11948 5972 12412
rect 6028 12403 6068 12412
rect 6315 12452 6357 12461
rect 8716 12452 8756 12461
rect 6315 12412 6316 12452
rect 6356 12412 6357 12452
rect 6315 12403 6357 12412
rect 8524 12412 8716 12452
rect 5932 11899 5972 11908
rect 6124 11780 6164 11789
rect 6124 11360 6164 11740
rect 5836 11320 6164 11360
rect 6316 11360 6356 12403
rect 6412 12284 6452 12293
rect 6412 11780 6452 12244
rect 7276 12284 7316 12293
rect 6508 11780 6548 11789
rect 6412 11740 6508 11780
rect 6508 11731 6548 11740
rect 7276 11360 7316 12244
rect 8524 11948 8564 12412
rect 8716 12403 8756 12412
rect 9388 12284 9428 12293
rect 9428 12244 9524 12284
rect 9388 12235 9428 12244
rect 8524 11899 8564 11908
rect 6316 11320 6452 11360
rect 5836 11024 5876 11320
rect 5836 10975 5876 10984
rect 5452 10891 5492 10900
rect 5548 10940 5588 10949
rect 5068 10772 5108 10781
rect 5108 10732 5396 10772
rect 5068 10723 5108 10732
rect 4779 10604 4821 10613
rect 4779 10564 4780 10604
rect 4820 10564 4821 10604
rect 4779 10555 4821 10564
rect 4928 10604 5296 10613
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 4928 10555 5296 10564
rect 4876 10436 4916 10445
rect 4684 10396 4876 10436
rect 4876 10387 4916 10396
rect 5067 10436 5109 10445
rect 5356 10436 5396 10732
rect 5548 10436 5588 10900
rect 6412 10940 6452 11320
rect 6412 10891 6452 10900
rect 7180 11320 7316 11360
rect 7372 11780 7412 11789
rect 6892 10772 6932 10781
rect 5067 10396 5068 10436
rect 5108 10396 5109 10436
rect 5067 10387 5109 10396
rect 5164 10396 5396 10436
rect 5452 10396 5588 10436
rect 5836 10436 5876 10445
rect 5876 10396 6260 10436
rect 5068 10302 5108 10387
rect 4395 10268 4437 10277
rect 4395 10228 4396 10268
rect 4436 10228 4437 10268
rect 4395 10219 4437 10228
rect 5164 10268 5204 10396
rect 5164 10219 5204 10228
rect 5260 10268 5300 10277
rect 4396 9680 4436 10219
rect 5260 10109 5300 10228
rect 5355 10268 5397 10277
rect 5452 10268 5492 10396
rect 5836 10387 5876 10396
rect 5355 10228 5356 10268
rect 5396 10228 5492 10268
rect 5548 10268 5588 10277
rect 5355 10219 5397 10228
rect 5356 10134 5396 10219
rect 5259 10100 5301 10109
rect 5259 10060 5260 10100
rect 5300 10060 5301 10100
rect 5259 10051 5301 10060
rect 4396 9631 4436 9640
rect 4491 9512 4533 9521
rect 4491 9472 4492 9512
rect 4532 9472 4533 9512
rect 4491 9463 4533 9472
rect 4300 9379 4340 9388
rect 4492 9428 4532 9463
rect 4492 8933 4532 9388
rect 4683 9428 4725 9437
rect 4683 9388 4684 9428
rect 4724 9388 4725 9428
rect 4683 9379 4725 9388
rect 5068 9428 5108 9437
rect 5548 9428 5588 10228
rect 5644 10268 5684 10277
rect 5644 9605 5684 10228
rect 5740 10268 5780 10277
rect 5643 9596 5685 9605
rect 5643 9556 5644 9596
rect 5684 9556 5685 9596
rect 5643 9547 5685 9556
rect 5108 9388 5396 9428
rect 5548 9388 5684 9428
rect 5068 9379 5108 9388
rect 4684 9294 4724 9379
rect 5164 9260 5204 9269
rect 4780 9220 5164 9260
rect 4491 8924 4533 8933
rect 4108 8884 4244 8924
rect 3243 8840 3285 8849
rect 3628 8840 3668 8849
rect 3243 8800 3244 8840
rect 3284 8800 3285 8840
rect 3243 8791 3285 8800
rect 3532 8800 3628 8840
rect 2612 7876 2708 7916
rect 2572 7867 2612 7876
rect 2956 7832 2996 8716
rect 3148 8707 3188 8716
rect 3244 8706 3284 8791
rect 3340 8756 3380 8767
rect 3340 8681 3380 8716
rect 3339 8672 3381 8681
rect 3339 8632 3340 8672
rect 3380 8632 3381 8672
rect 3339 8623 3381 8632
rect 2668 7792 2996 7832
rect 3436 7916 3476 7925
rect 1419 7748 1461 7757
rect 1419 7708 1420 7748
rect 1460 7708 1461 7748
rect 1419 7699 1461 7708
rect 1899 7748 1941 7757
rect 1899 7708 1900 7748
rect 1940 7708 1941 7748
rect 1899 7699 1941 7708
rect 1420 7244 1460 7699
rect 1516 7244 1556 7253
rect 1420 7204 1516 7244
rect 1131 6992 1173 7001
rect 1131 6952 1132 6992
rect 1172 6952 1173 6992
rect 1131 6943 1173 6952
rect 1132 5648 1172 6943
rect 1227 6404 1269 6413
rect 1227 6364 1228 6404
rect 1268 6364 1269 6404
rect 1227 6355 1269 6364
rect 1228 6270 1268 6355
rect 1324 5741 1364 7204
rect 1516 7195 1556 7204
rect 1708 7244 1748 7253
rect 1611 7160 1653 7169
rect 1611 7120 1612 7160
rect 1652 7120 1653 7160
rect 1611 7111 1653 7120
rect 1612 7026 1652 7111
rect 1708 7085 1748 7204
rect 1900 7244 1940 7699
rect 1995 7328 2037 7337
rect 1995 7288 1996 7328
rect 2036 7288 2037 7328
rect 1995 7279 2037 7288
rect 1900 7195 1940 7204
rect 1996 7194 2036 7279
rect 2092 7244 2132 7253
rect 2092 7085 2132 7204
rect 1707 7076 1749 7085
rect 1707 7036 1708 7076
rect 1748 7036 1749 7076
rect 1707 7027 1749 7036
rect 2091 7076 2133 7085
rect 2091 7036 2092 7076
rect 2132 7036 2133 7076
rect 2091 7027 2133 7036
rect 2284 6992 2324 7001
rect 2284 6413 2324 6952
rect 1612 6404 1652 6413
rect 2283 6404 2325 6413
rect 1652 6364 1748 6404
rect 1612 6355 1652 6364
rect 1419 5984 1461 5993
rect 1419 5944 1420 5984
rect 1460 5944 1461 5984
rect 1419 5935 1461 5944
rect 1420 5900 1460 5935
rect 1420 5849 1460 5860
rect 1611 5816 1653 5825
rect 1611 5776 1612 5816
rect 1652 5776 1653 5816
rect 1611 5767 1653 5776
rect 1323 5732 1365 5741
rect 1323 5692 1324 5732
rect 1364 5692 1365 5732
rect 1323 5683 1365 5692
rect 1228 5648 1268 5657
rect 1132 5608 1228 5648
rect 1228 5599 1268 5608
rect 1612 5648 1652 5767
rect 1708 5732 1748 6364
rect 2283 6364 2284 6404
rect 2324 6364 2325 6404
rect 2283 6355 2325 6364
rect 2475 6404 2517 6413
rect 2475 6364 2476 6404
rect 2516 6364 2517 6404
rect 2475 6355 2517 6364
rect 2476 6270 2516 6355
rect 1804 5900 1844 5909
rect 1844 5860 2516 5900
rect 1804 5851 1844 5860
rect 1996 5732 2036 5741
rect 1708 5692 1996 5732
rect 1996 5683 2036 5692
rect 2091 5732 2133 5741
rect 2091 5692 2092 5732
rect 2132 5692 2133 5732
rect 2091 5683 2133 5692
rect 2476 5732 2516 5860
rect 2476 5683 2516 5692
rect 2571 5732 2613 5741
rect 2571 5692 2572 5732
rect 2612 5692 2613 5732
rect 2571 5683 2613 5692
rect 2668 5732 2708 7792
rect 3436 7589 3476 7876
rect 3435 7580 3477 7589
rect 3435 7540 3436 7580
rect 3476 7540 3477 7580
rect 3435 7531 3477 7540
rect 3436 7412 3476 7421
rect 2956 7372 3436 7412
rect 2956 7244 2996 7372
rect 3436 7363 3476 7372
rect 2956 7195 2996 7204
rect 3148 7244 3188 7253
rect 2859 5816 2901 5825
rect 2859 5776 2860 5816
rect 2900 5776 2901 5816
rect 2859 5767 2901 5776
rect 2668 5683 2708 5692
rect 2860 5732 2900 5767
rect 3148 5741 3188 7204
rect 3244 7244 3284 7253
rect 3244 7085 3284 7204
rect 3339 7244 3381 7253
rect 3339 7204 3340 7244
rect 3380 7204 3381 7244
rect 3339 7195 3381 7204
rect 3340 7110 3380 7195
rect 3243 7076 3285 7085
rect 3243 7036 3244 7076
rect 3284 7036 3285 7076
rect 3243 7027 3285 7036
rect 3532 6824 3572 8800
rect 3628 8791 3668 8800
rect 3820 8756 3860 8765
rect 3820 8504 3860 8716
rect 4107 8756 4149 8765
rect 4107 8716 4108 8756
rect 4148 8716 4149 8756
rect 4107 8707 4149 8716
rect 4108 8622 4148 8707
rect 3820 8464 4148 8504
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 4012 8168 4052 8177
rect 4108 8168 4148 8464
rect 4052 8128 4148 8168
rect 4012 8119 4052 8128
rect 4204 7925 4244 8884
rect 4491 8884 4492 8924
rect 4532 8884 4533 8924
rect 4491 8875 4533 8884
rect 4300 8756 4340 8765
rect 4300 8597 4340 8716
rect 4491 8756 4533 8765
rect 4491 8716 4492 8756
rect 4532 8716 4533 8756
rect 4491 8707 4533 8716
rect 4588 8756 4628 8767
rect 4299 8588 4341 8597
rect 4299 8548 4300 8588
rect 4340 8548 4341 8588
rect 4299 8539 4341 8548
rect 4396 8504 4436 8513
rect 4203 7916 4245 7925
rect 4203 7876 4204 7916
rect 4244 7876 4245 7916
rect 4203 7867 4245 7876
rect 3820 7832 3860 7841
rect 3820 7421 3860 7792
rect 4299 7664 4341 7673
rect 4299 7624 4300 7664
rect 4340 7624 4341 7664
rect 4299 7615 4341 7624
rect 3819 7412 3861 7421
rect 3819 7372 3820 7412
rect 3860 7372 3861 7412
rect 3819 7363 3861 7372
rect 3819 7244 3861 7253
rect 3819 7204 3820 7244
rect 3860 7204 3861 7244
rect 3819 7195 3861 7204
rect 3820 7110 3860 7195
rect 3436 6784 3572 6824
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 1612 5599 1652 5608
rect 2092 5598 2132 5683
rect 2572 5598 2612 5683
rect 2764 4892 2804 4901
rect 2860 4892 2900 5692
rect 3052 5732 3092 5741
rect 2955 5648 2997 5657
rect 2955 5608 2956 5648
rect 2996 5608 2997 5648
rect 2955 5599 2997 5608
rect 2956 5514 2996 5599
rect 3052 4901 3092 5692
rect 3147 5732 3189 5741
rect 3147 5692 3148 5732
rect 3188 5692 3189 5732
rect 3147 5683 3189 5692
rect 3436 5732 3476 6784
rect 3688 6775 4056 6784
rect 3628 6488 3668 6497
rect 3668 6448 3860 6488
rect 3628 6439 3668 6448
rect 3820 6404 3860 6448
rect 3820 6355 3860 6364
rect 4300 5993 4340 7615
rect 4396 7589 4436 8464
rect 4395 7580 4437 7589
rect 4395 7540 4396 7580
rect 4436 7540 4437 7580
rect 4395 7531 4437 7540
rect 4492 7412 4532 8707
rect 4588 8681 4628 8716
rect 4587 8672 4629 8681
rect 4587 8632 4588 8672
rect 4628 8632 4629 8672
rect 4587 8623 4629 8632
rect 4587 7916 4629 7925
rect 4587 7876 4588 7916
rect 4628 7876 4629 7916
rect 4587 7867 4629 7876
rect 4684 7916 4724 7925
rect 4396 7372 4532 7412
rect 4396 7001 4436 7372
rect 4491 7244 4533 7253
rect 4491 7204 4492 7244
rect 4532 7204 4533 7244
rect 4491 7195 4533 7204
rect 4492 7110 4532 7195
rect 4395 6992 4437 7001
rect 4395 6952 4396 6992
rect 4436 6952 4437 6992
rect 4395 6943 4437 6952
rect 4396 6656 4436 6943
rect 4492 6656 4532 6665
rect 4396 6616 4492 6656
rect 4492 6607 4532 6616
rect 4299 5984 4341 5993
rect 4299 5944 4300 5984
rect 4340 5944 4341 5984
rect 4299 5935 4341 5944
rect 3819 5900 3861 5909
rect 3819 5860 3820 5900
rect 3860 5860 3861 5900
rect 3819 5851 3861 5860
rect 3820 5766 3860 5851
rect 4588 5741 4628 7867
rect 4684 7757 4724 7876
rect 4683 7748 4725 7757
rect 4683 7708 4684 7748
rect 4724 7708 4725 7748
rect 4683 7699 4725 7708
rect 4683 7412 4725 7421
rect 4683 7372 4684 7412
rect 4724 7372 4725 7412
rect 4683 7363 4725 7372
rect 4684 7278 4724 7363
rect 4780 7244 4820 9220
rect 5164 9211 5204 9220
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 5067 8924 5109 8933
rect 5067 8884 5068 8924
rect 5108 8884 5109 8924
rect 5067 8875 5109 8884
rect 5260 8924 5300 8933
rect 5356 8924 5396 9388
rect 5300 8884 5396 8924
rect 5548 9260 5588 9269
rect 5260 8875 5300 8884
rect 4971 8336 5013 8345
rect 4971 8296 4972 8336
rect 5012 8296 5013 8336
rect 4971 8287 5013 8296
rect 4972 8168 5012 8287
rect 4972 8119 5012 8128
rect 4876 7916 4916 7925
rect 4876 7757 4916 7876
rect 5068 7916 5108 8875
rect 5452 8840 5492 8849
rect 5548 8840 5588 9220
rect 5492 8800 5588 8840
rect 5452 8791 5492 8800
rect 5451 8588 5493 8597
rect 5451 8548 5452 8588
rect 5492 8548 5493 8588
rect 5451 8539 5493 8548
rect 5068 7867 5108 7876
rect 5260 7916 5300 7927
rect 5260 7841 5300 7876
rect 5259 7832 5301 7841
rect 5259 7792 5260 7832
rect 5300 7792 5301 7832
rect 5259 7783 5301 7792
rect 4875 7748 4917 7757
rect 4875 7708 4876 7748
rect 4916 7708 4917 7748
rect 4875 7699 4917 7708
rect 5356 7748 5396 7757
rect 5356 7589 5396 7708
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 5355 7580 5397 7589
rect 5355 7540 5356 7580
rect 5396 7540 5397 7580
rect 5355 7531 5397 7540
rect 5067 7412 5109 7421
rect 5067 7372 5068 7412
rect 5108 7372 5109 7412
rect 5067 7363 5109 7372
rect 4876 7244 4916 7253
rect 4780 7204 4876 7244
rect 4876 7195 4916 7204
rect 4971 7244 5013 7253
rect 4971 7204 4972 7244
rect 5012 7204 5013 7244
rect 4971 7195 5013 7204
rect 4972 7110 5012 7195
rect 4779 6404 4821 6413
rect 4779 6364 4780 6404
rect 4820 6364 4821 6404
rect 4779 6355 4821 6364
rect 5068 6404 5108 7363
rect 5452 7244 5492 8539
rect 5644 8345 5684 9388
rect 5643 8336 5685 8345
rect 5643 8296 5644 8336
rect 5684 8296 5685 8336
rect 5643 8287 5685 8296
rect 5548 8168 5588 8177
rect 5740 8168 5780 10228
rect 6123 10268 6165 10277
rect 6123 10228 6124 10268
rect 6164 10228 6165 10268
rect 6123 10219 6165 10228
rect 6028 10016 6068 10025
rect 5836 9976 6028 10016
rect 5836 8756 5876 9976
rect 6028 9967 6068 9976
rect 5931 9596 5973 9605
rect 5931 9556 5932 9596
rect 5972 9556 5973 9596
rect 5931 9547 5973 9556
rect 5932 8849 5972 9547
rect 5931 8840 5973 8849
rect 5931 8800 5932 8840
rect 5972 8800 5973 8840
rect 5931 8791 5973 8800
rect 5836 8707 5876 8716
rect 6124 8597 6164 10219
rect 6220 9428 6260 10396
rect 6892 10277 6932 10732
rect 6891 10268 6933 10277
rect 6891 10228 6892 10268
rect 6932 10228 6933 10268
rect 6891 10219 6933 10228
rect 6988 10268 7028 10277
rect 6699 10100 6741 10109
rect 6699 10060 6700 10100
rect 6740 10060 6741 10100
rect 6699 10051 6741 10060
rect 6220 9379 6260 9388
rect 6411 9428 6453 9437
rect 6411 9388 6412 9428
rect 6452 9388 6453 9428
rect 6411 9379 6453 9388
rect 6604 9428 6644 9437
rect 6412 9294 6452 9379
rect 6508 9344 6548 9353
rect 6123 8588 6165 8597
rect 6508 8588 6548 9304
rect 6604 8681 6644 9388
rect 6700 8756 6740 10051
rect 6988 9521 7028 10228
rect 7180 10268 7220 11320
rect 7180 10219 7220 10228
rect 7083 10184 7125 10193
rect 7083 10144 7084 10184
rect 7124 10144 7125 10184
rect 7083 10135 7125 10144
rect 7084 10050 7124 10135
rect 7372 10109 7412 11740
rect 8235 11780 8277 11789
rect 8235 11740 8236 11780
rect 8276 11740 8277 11780
rect 8235 11731 8277 11740
rect 9388 11780 9428 11789
rect 9484 11780 9524 12244
rect 9580 11789 9620 11874
rect 9579 11780 9621 11789
rect 9484 11740 9580 11780
rect 9620 11740 9621 11780
rect 7563 11696 7605 11705
rect 7563 11656 7564 11696
rect 7604 11656 7605 11696
rect 7563 11647 7605 11656
rect 7564 10940 7604 11647
rect 7564 10891 7604 10900
rect 7756 10940 7796 10949
rect 8236 10940 8276 11731
rect 9388 11612 9428 11740
rect 9579 11731 9621 11740
rect 9772 11780 9812 11791
rect 9772 11705 9812 11740
rect 10636 11780 10676 11791
rect 10636 11705 10676 11740
rect 9771 11696 9813 11705
rect 9771 11656 9772 11696
rect 9812 11656 9813 11696
rect 9771 11647 9813 11656
rect 10635 11696 10677 11705
rect 10635 11656 10636 11696
rect 10676 11656 10677 11696
rect 10635 11647 10677 11656
rect 11115 11696 11157 11705
rect 11115 11656 11116 11696
rect 11156 11656 11157 11696
rect 11115 11647 11157 11656
rect 9676 11612 9716 11621
rect 9388 11572 9676 11612
rect 9676 11563 9716 11572
rect 8523 11528 8565 11537
rect 8523 11488 8524 11528
rect 8564 11488 8565 11528
rect 8523 11479 8565 11488
rect 8716 11528 8756 11537
rect 7796 10900 8236 10940
rect 7756 10891 7796 10900
rect 8236 10891 8276 10900
rect 8524 10940 8564 11479
rect 8716 11360 8756 11488
rect 9963 11528 10005 11537
rect 9963 11488 9964 11528
rect 10004 11488 10005 11528
rect 9963 11479 10005 11488
rect 9964 11394 10004 11479
rect 8524 10891 8564 10900
rect 8620 11320 8756 11360
rect 7660 10772 7700 10781
rect 8044 10772 8084 10781
rect 8620 10772 8660 11320
rect 11116 11192 11156 11647
rect 11116 11143 11156 11152
rect 9100 10940 9140 10949
rect 7660 10445 7700 10732
rect 7756 10732 8044 10772
rect 7659 10436 7701 10445
rect 7659 10396 7660 10436
rect 7700 10396 7701 10436
rect 7659 10387 7701 10396
rect 7660 10268 7700 10277
rect 7660 10193 7700 10228
rect 7756 10268 7796 10732
rect 8044 10723 8084 10732
rect 8524 10732 8660 10772
rect 8716 10856 8756 10865
rect 8043 10436 8085 10445
rect 8043 10396 8044 10436
rect 8084 10396 8085 10436
rect 8043 10387 8085 10396
rect 7756 10219 7796 10228
rect 7659 10184 7701 10193
rect 7659 10144 7660 10184
rect 7700 10144 7701 10184
rect 7659 10135 7701 10144
rect 7948 10184 7988 10193
rect 7371 10100 7413 10109
rect 7371 10060 7372 10100
rect 7412 10060 7413 10100
rect 7371 10051 7413 10060
rect 7660 9941 7700 10135
rect 7659 9932 7701 9941
rect 7659 9892 7660 9932
rect 7700 9892 7701 9932
rect 7659 9883 7701 9892
rect 6987 9512 7029 9521
rect 6987 9472 6988 9512
rect 7028 9472 7029 9512
rect 6987 9463 7029 9472
rect 6795 9428 6837 9437
rect 6795 9388 6796 9428
rect 6836 9388 6837 9428
rect 6795 9379 6837 9388
rect 6796 9294 6836 9379
rect 6700 8707 6740 8716
rect 6603 8672 6645 8681
rect 6603 8632 6604 8672
rect 6644 8632 6645 8672
rect 6603 8623 6645 8632
rect 6123 8548 6124 8588
rect 6164 8548 6165 8588
rect 6123 8539 6165 8548
rect 6220 8548 6548 8588
rect 5588 8128 5780 8168
rect 5548 8119 5588 8128
rect 6220 7916 6260 8548
rect 6220 7867 6260 7876
rect 6411 7916 6453 7925
rect 6411 7876 6412 7916
rect 6452 7876 6453 7916
rect 6411 7867 6453 7876
rect 5835 7832 5877 7841
rect 5835 7792 5836 7832
rect 5876 7792 5877 7832
rect 5835 7783 5877 7792
rect 5548 7244 5588 7253
rect 5452 7204 5548 7244
rect 5548 7195 5588 7204
rect 5836 7076 5876 7783
rect 6412 7782 6452 7867
rect 6604 7412 6644 8623
rect 6988 8597 7028 9463
rect 7948 9437 7988 10144
rect 8044 10100 8084 10387
rect 8140 10268 8180 10277
rect 8180 10228 8468 10268
rect 8140 10219 8180 10228
rect 8044 10060 8276 10100
rect 8139 9932 8181 9941
rect 8139 9892 8140 9932
rect 8180 9892 8181 9932
rect 8139 9883 8181 9892
rect 7468 9428 7508 9437
rect 7468 8849 7508 9388
rect 7852 9428 7892 9437
rect 7852 9008 7892 9388
rect 7947 9428 7989 9437
rect 7947 9388 7948 9428
rect 7988 9388 7989 9428
rect 7947 9379 7989 9388
rect 8140 9428 8180 9883
rect 8140 9379 8180 9388
rect 8236 9428 8276 10060
rect 8236 9379 8276 9388
rect 8332 9428 8372 9437
rect 7947 9260 7989 9269
rect 7947 9220 7948 9260
rect 7988 9220 7989 9260
rect 8332 9260 8372 9388
rect 8428 9428 8468 10228
rect 8428 9379 8468 9388
rect 8524 9260 8564 10732
rect 8716 10436 8756 10816
rect 8812 10436 8852 10445
rect 8716 10396 8812 10436
rect 8812 10387 8852 10396
rect 8619 9428 8661 9437
rect 8619 9388 8620 9428
rect 8660 9388 8661 9428
rect 8619 9379 8661 9388
rect 9004 9428 9044 9437
rect 8620 9294 8660 9379
rect 9004 9269 9044 9388
rect 8332 9220 8564 9260
rect 9003 9260 9045 9269
rect 9003 9220 9004 9260
rect 9044 9220 9045 9260
rect 7947 9211 7989 9220
rect 9003 9211 9045 9220
rect 7948 9126 7988 9211
rect 9100 9008 9140 10900
rect 9964 10940 10004 10949
rect 9964 10352 10004 10900
rect 9964 10303 10004 10312
rect 10252 10396 10676 10436
rect 7852 8968 7988 9008
rect 7467 8840 7509 8849
rect 7467 8800 7468 8840
rect 7508 8800 7509 8840
rect 7467 8791 7509 8800
rect 7851 8840 7893 8849
rect 7851 8800 7852 8840
rect 7892 8800 7893 8840
rect 7851 8791 7893 8800
rect 7852 8672 7892 8791
rect 7852 8623 7892 8632
rect 6987 8588 7029 8597
rect 6987 8548 6988 8588
rect 7028 8548 7029 8588
rect 6987 8539 7029 8548
rect 7563 8588 7605 8597
rect 7563 8548 7564 8588
rect 7604 8548 7605 8588
rect 7563 8539 7605 8548
rect 7083 8168 7125 8177
rect 7083 8128 7084 8168
rect 7124 8128 7125 8168
rect 7083 8119 7125 8128
rect 7084 8034 7124 8119
rect 7276 7916 7316 7925
rect 6796 7412 6836 7421
rect 6604 7372 6796 7412
rect 6796 7363 6836 7372
rect 5836 7027 5876 7036
rect 6220 6992 6260 7001
rect 5068 6355 5108 6364
rect 5931 6404 5973 6413
rect 5931 6364 5932 6404
rect 5972 6364 5973 6404
rect 5931 6355 5973 6364
rect 4684 6320 4724 6329
rect 4684 5909 4724 6280
rect 4683 5900 4725 5909
rect 4683 5860 4684 5900
rect 4724 5860 4725 5900
rect 4683 5851 4725 5860
rect 3436 5683 3476 5692
rect 3531 5732 3573 5741
rect 3531 5692 3532 5732
rect 3572 5692 3573 5732
rect 3531 5683 3573 5692
rect 4587 5732 4629 5741
rect 4587 5692 4588 5732
rect 4628 5692 4629 5732
rect 4587 5683 4629 5692
rect 3532 5598 3572 5683
rect 4684 5480 4724 5489
rect 4780 5480 4820 6355
rect 5643 6320 5685 6329
rect 5643 6280 5644 6320
rect 5684 6280 5685 6320
rect 5643 6271 5685 6280
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 4875 5732 4917 5741
rect 4875 5692 4876 5732
rect 4916 5692 4917 5732
rect 4875 5683 4917 5692
rect 4876 5598 4916 5683
rect 4724 5440 4820 5480
rect 5260 5480 5300 5489
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 3339 5060 3381 5069
rect 3339 5020 3340 5060
rect 3380 5020 3381 5060
rect 3339 5011 3381 5020
rect 3147 4976 3189 4985
rect 3147 4936 3148 4976
rect 3188 4936 3189 4976
rect 3147 4927 3189 4936
rect 2804 4852 2900 4892
rect 2956 4892 2996 4901
rect 3051 4892 3093 4901
rect 2996 4852 3052 4892
rect 3092 4852 3093 4892
rect 2764 4843 2804 4852
rect 2956 4843 2996 4852
rect 3051 4843 3093 4852
rect 3148 4892 3188 4927
rect 3148 4841 3188 4852
rect 3244 4892 3284 4901
rect 2860 4724 2900 4733
rect 3244 4724 3284 4852
rect 3340 4892 3380 5011
rect 3340 4843 3380 4852
rect 3435 4892 3477 4901
rect 3435 4852 3436 4892
rect 3476 4852 3477 4892
rect 3435 4843 3477 4852
rect 4299 4892 4341 4901
rect 4299 4852 4300 4892
rect 4340 4852 4341 4892
rect 4299 4843 4341 4852
rect 4587 4892 4629 4901
rect 4587 4852 4588 4892
rect 4628 4852 4629 4892
rect 4587 4843 4629 4852
rect 3436 4758 3476 4843
rect 4300 4758 4340 4843
rect 3628 4724 3668 4733
rect 2900 4684 3284 4724
rect 3532 4684 3628 4724
rect 2860 4675 2900 4684
rect 3532 4472 3572 4684
rect 3628 4675 3668 4684
rect 2668 4432 3572 4472
rect 2668 4304 2708 4432
rect 2668 4255 2708 4264
rect 3052 4220 3092 4229
rect 3052 3632 3092 4180
rect 3916 4220 3956 4229
rect 3916 4061 3956 4180
rect 4588 4145 4628 4843
rect 4587 4136 4629 4145
rect 4587 4096 4588 4136
rect 4628 4096 4629 4136
rect 4587 4087 4629 4096
rect 4684 4061 4724 5440
rect 5260 5069 5300 5440
rect 5451 5480 5493 5489
rect 5451 5440 5452 5480
rect 5492 5440 5493 5480
rect 5451 5431 5493 5440
rect 5259 5060 5301 5069
rect 5259 5020 5260 5060
rect 5300 5020 5301 5060
rect 5259 5011 5301 5020
rect 4780 4901 4820 4986
rect 4779 4892 4821 4901
rect 4779 4852 4780 4892
rect 4820 4852 4821 4892
rect 4779 4843 4821 4852
rect 4876 4892 4916 4901
rect 4876 4724 4916 4852
rect 5260 4892 5300 4901
rect 5300 4852 5396 4892
rect 5260 4843 5300 4852
rect 5068 4733 5108 4818
rect 4780 4684 4916 4724
rect 5067 4724 5109 4733
rect 5067 4684 5068 4724
rect 5108 4684 5109 4724
rect 4780 4313 4820 4684
rect 5067 4675 5109 4684
rect 5356 4565 5396 4852
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 5355 4556 5397 4565
rect 5355 4516 5356 4556
rect 5396 4516 5397 4556
rect 5355 4507 5397 4516
rect 5067 4388 5109 4397
rect 5067 4348 5068 4388
rect 5108 4348 5109 4388
rect 5067 4339 5109 4348
rect 4779 4304 4821 4313
rect 4779 4264 4780 4304
rect 4820 4264 4821 4304
rect 4779 4255 4821 4264
rect 5068 4254 5108 4339
rect 5259 4304 5301 4313
rect 5356 4304 5396 4313
rect 5259 4264 5260 4304
rect 5300 4264 5356 4304
rect 5259 4255 5301 4264
rect 5356 4255 5396 4264
rect 5452 4220 5492 5431
rect 5547 4724 5589 4733
rect 5547 4684 5548 4724
rect 5588 4684 5589 4724
rect 5547 4675 5589 4684
rect 5452 4171 5492 4180
rect 5163 4136 5205 4145
rect 5163 4096 5164 4136
rect 5204 4096 5205 4136
rect 5163 4087 5205 4096
rect 3915 4052 3957 4061
rect 3915 4012 3916 4052
rect 3956 4012 3957 4052
rect 3915 4003 3957 4012
rect 4683 4052 4725 4061
rect 4683 4012 4684 4052
rect 4724 4012 4725 4052
rect 4683 4003 4725 4012
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 3243 3716 3285 3725
rect 3243 3676 3244 3716
rect 3284 3676 3285 3716
rect 3243 3667 3285 3676
rect 3148 3632 3188 3641
rect 3052 3592 3148 3632
rect 3148 3583 3188 3592
rect 3244 3380 3284 3667
rect 5164 3632 5204 4087
rect 5164 3583 5204 3592
rect 5067 3464 5109 3473
rect 5067 3424 5068 3464
rect 5108 3424 5109 3464
rect 5067 3415 5109 3424
rect 3244 3331 3284 3340
rect 5068 3380 5108 3415
rect 5068 3329 5108 3340
rect 5259 3380 5301 3389
rect 5259 3340 5260 3380
rect 5300 3340 5301 3380
rect 5259 3331 5301 3340
rect 5452 3380 5492 3389
rect 5548 3380 5588 4675
rect 5644 3473 5684 6271
rect 5932 6270 5972 6355
rect 5932 5732 5972 5743
rect 5932 5657 5972 5692
rect 6220 5732 6260 6952
rect 7084 6236 7124 6245
rect 6891 5900 6933 5909
rect 6891 5860 6892 5900
rect 6932 5860 6933 5900
rect 6891 5851 6933 5860
rect 6220 5657 6260 5692
rect 6603 5732 6645 5741
rect 6603 5692 6604 5732
rect 6644 5692 6645 5732
rect 6603 5683 6645 5692
rect 5931 5648 5973 5657
rect 5931 5608 5932 5648
rect 5972 5608 5973 5648
rect 5931 5599 5973 5608
rect 6219 5648 6261 5657
rect 6219 5608 6220 5648
rect 6260 5608 6261 5648
rect 6219 5599 6261 5608
rect 6124 5480 6164 5489
rect 6028 5440 6124 5480
rect 5931 4808 5973 4817
rect 5836 4768 5932 4808
rect 5972 4768 5973 4808
rect 5836 4220 5876 4768
rect 5931 4759 5973 4768
rect 5932 4674 5972 4759
rect 5836 4171 5876 4180
rect 5643 3464 5685 3473
rect 5643 3424 5644 3464
rect 5684 3424 5685 3464
rect 5643 3415 5685 3424
rect 5492 3340 5588 3380
rect 5836 3380 5876 3389
rect 6028 3380 6068 5440
rect 6124 5431 6164 5440
rect 6124 4892 6164 4901
rect 6220 4892 6260 5599
rect 6411 5480 6453 5489
rect 6411 5440 6412 5480
rect 6452 5440 6453 5480
rect 6411 5431 6453 5440
rect 6412 5346 6452 5431
rect 6411 5060 6453 5069
rect 6411 5020 6412 5060
rect 6452 5020 6453 5060
rect 6411 5011 6453 5020
rect 6164 4852 6260 4892
rect 6412 4892 6452 5011
rect 6124 3725 6164 4852
rect 6219 4724 6261 4733
rect 6219 4684 6220 4724
rect 6260 4684 6261 4724
rect 6219 4675 6261 4684
rect 6220 4590 6260 4675
rect 6315 4388 6357 4397
rect 6315 4348 6316 4388
rect 6356 4348 6357 4388
rect 6315 4339 6357 4348
rect 6316 4304 6356 4339
rect 6316 4253 6356 4264
rect 6220 4220 6260 4229
rect 6220 3809 6260 4180
rect 6412 4220 6452 4852
rect 6604 4388 6644 5683
rect 6795 5480 6837 5489
rect 6795 5440 6796 5480
rect 6836 5440 6837 5480
rect 6795 5431 6837 5440
rect 6699 4892 6741 4901
rect 6699 4852 6700 4892
rect 6740 4852 6741 4892
rect 6699 4843 6741 4852
rect 6700 4758 6740 4843
rect 6699 4472 6741 4481
rect 6699 4432 6700 4472
rect 6740 4432 6741 4472
rect 6699 4423 6741 4432
rect 6604 4339 6644 4348
rect 6412 4171 6452 4180
rect 6700 4220 6740 4423
rect 6700 4171 6740 4180
rect 6796 4220 6836 5431
rect 6892 4808 6932 5851
rect 7084 5825 7124 6196
rect 7276 6152 7316 7876
rect 7564 7580 7604 8539
rect 7948 8168 7988 8968
rect 8812 8968 9140 9008
rect 9196 10268 9236 10277
rect 8812 8924 8852 8968
rect 8716 8884 8852 8924
rect 8620 8840 8660 8849
rect 8716 8840 8756 8884
rect 8660 8800 8756 8840
rect 8907 8840 8949 8849
rect 8907 8800 8908 8840
rect 8948 8800 8949 8840
rect 8620 8791 8660 8800
rect 8907 8791 8949 8800
rect 8236 8756 8276 8765
rect 8524 8756 8564 8765
rect 8812 8756 8852 8765
rect 8276 8716 8524 8756
rect 8236 8168 8276 8716
rect 8524 8707 8564 8716
rect 8716 8716 8812 8756
rect 8427 8588 8469 8597
rect 8427 8548 8428 8588
rect 8468 8548 8469 8588
rect 8427 8539 8469 8548
rect 7372 7540 7604 7580
rect 7852 8128 8276 8168
rect 8332 8504 8372 8513
rect 7372 6404 7412 7540
rect 7372 6329 7412 6364
rect 7563 6404 7605 6413
rect 7563 6364 7564 6404
rect 7604 6364 7605 6404
rect 7563 6355 7605 6364
rect 7371 6320 7413 6329
rect 7371 6280 7372 6320
rect 7412 6280 7413 6320
rect 7371 6271 7413 6280
rect 7468 6320 7508 6329
rect 7372 6240 7412 6271
rect 7468 6245 7508 6280
rect 7564 6270 7604 6355
rect 7467 6236 7509 6245
rect 7467 6196 7468 6236
rect 7508 6196 7509 6236
rect 7467 6187 7509 6196
rect 7276 6112 7412 6152
rect 7083 5816 7125 5825
rect 7083 5776 7084 5816
rect 7124 5776 7125 5816
rect 7083 5767 7125 5776
rect 7084 5732 7124 5767
rect 7084 5682 7124 5692
rect 7083 5564 7125 5573
rect 7083 5524 7084 5564
rect 7124 5524 7125 5564
rect 7083 5515 7125 5524
rect 6892 4759 6932 4768
rect 7084 4388 7124 5515
rect 7276 5480 7316 5489
rect 7180 4724 7220 4733
rect 7180 4481 7220 4684
rect 7179 4472 7221 4481
rect 7179 4432 7180 4472
rect 7220 4432 7221 4472
rect 7179 4423 7221 4432
rect 6796 4171 6836 4180
rect 6892 4348 7124 4388
rect 6892 4220 6932 4348
rect 6892 4171 6932 4180
rect 7084 4220 7124 4229
rect 7276 4220 7316 5440
rect 7372 4313 7412 6112
rect 7468 5573 7508 6187
rect 7852 5657 7892 8128
rect 7947 8000 7989 8009
rect 7947 7960 7948 8000
rect 7988 7960 7989 8000
rect 7947 7951 7989 7960
rect 7948 7916 7988 7951
rect 8332 7925 8372 8464
rect 7948 7865 7988 7876
rect 8044 7916 8084 7925
rect 8044 7673 8084 7876
rect 8331 7916 8373 7925
rect 8331 7876 8332 7916
rect 8372 7876 8373 7916
rect 8331 7867 8373 7876
rect 8428 7916 8468 8539
rect 8524 8168 8564 8177
rect 8716 8168 8756 8716
rect 8812 8707 8852 8716
rect 8908 8756 8948 8791
rect 8908 8705 8948 8716
rect 9004 8756 9044 8767
rect 9004 8681 9044 8716
rect 9099 8756 9141 8765
rect 9099 8716 9100 8756
rect 9140 8716 9141 8756
rect 9099 8707 9141 8716
rect 9003 8672 9045 8681
rect 9003 8632 9004 8672
rect 9044 8632 9045 8672
rect 9003 8623 9045 8632
rect 9100 8622 9140 8707
rect 8907 8504 8949 8513
rect 8907 8464 8908 8504
rect 8948 8464 8949 8504
rect 8907 8455 8949 8464
rect 8564 8128 8756 8168
rect 8524 8009 8564 8128
rect 8523 8000 8565 8009
rect 8715 8000 8757 8009
rect 8523 7960 8524 8000
rect 8564 7960 8565 8000
rect 8523 7951 8565 7960
rect 8620 7960 8716 8000
rect 8756 7960 8757 8000
rect 8428 7867 8468 7876
rect 8620 7916 8660 7960
rect 8715 7951 8757 7960
rect 8620 7867 8660 7876
rect 8908 7916 8948 8455
rect 9196 8177 9236 10228
rect 10252 10268 10292 10396
rect 10252 10219 10292 10228
rect 10443 10268 10485 10277
rect 10443 10228 10444 10268
rect 10484 10228 10485 10268
rect 10443 10219 10485 10228
rect 10444 10134 10484 10219
rect 9387 10100 9429 10109
rect 9387 10060 9388 10100
rect 9428 10060 9429 10100
rect 9387 10051 9429 10060
rect 10636 10100 10676 10396
rect 11019 10268 11061 10277
rect 11019 10228 11020 10268
rect 11060 10228 11061 10268
rect 11019 10219 11061 10228
rect 11308 10268 11348 10277
rect 10676 10060 10964 10100
rect 10636 10051 10676 10060
rect 9388 9966 9428 10051
rect 9772 10016 9812 10025
rect 9772 9428 9812 9976
rect 10348 10016 10388 10025
rect 10388 9976 10580 10016
rect 10348 9967 10388 9976
rect 9868 9428 9908 9437
rect 9772 9388 9868 9428
rect 9868 9379 9908 9388
rect 9963 8756 10005 8765
rect 9963 8716 9964 8756
rect 10004 8716 10005 8756
rect 10540 8756 10580 9976
rect 10828 8756 10868 8765
rect 10540 8716 10828 8756
rect 9963 8707 10005 8716
rect 10828 8707 10868 8716
rect 9964 8622 10004 8707
rect 10155 8672 10197 8681
rect 10155 8632 10156 8672
rect 10196 8632 10197 8672
rect 10155 8623 10197 8632
rect 10156 8538 10196 8623
rect 10924 8588 10964 10060
rect 11020 9680 11060 10219
rect 11020 9631 11060 9640
rect 11020 9260 11060 9269
rect 11020 9008 11060 9220
rect 11020 8968 11252 9008
rect 11115 8840 11157 8849
rect 11115 8800 11116 8840
rect 11156 8800 11157 8840
rect 11115 8791 11157 8800
rect 11020 8756 11060 8765
rect 11020 8588 11060 8716
rect 11116 8706 11156 8791
rect 11212 8756 11252 8968
rect 10540 8548 11060 8588
rect 9291 8504 9333 8513
rect 9291 8464 9292 8504
rect 9332 8464 9333 8504
rect 9291 8455 9333 8464
rect 9292 8370 9332 8455
rect 9195 8168 9237 8177
rect 9195 8128 9196 8168
rect 9236 8128 9237 8168
rect 9195 8119 9237 8128
rect 9483 8168 9525 8177
rect 9483 8128 9484 8168
rect 9524 8128 9525 8168
rect 9483 8119 9525 8128
rect 8908 7867 8948 7876
rect 9291 7916 9333 7925
rect 9291 7876 9292 7916
rect 9332 7876 9333 7916
rect 9291 7867 9333 7876
rect 9292 7782 9332 7867
rect 8235 7748 8277 7757
rect 8235 7708 8236 7748
rect 8276 7708 8277 7748
rect 8235 7699 8277 7708
rect 9195 7748 9237 7757
rect 9195 7708 9196 7748
rect 9236 7708 9237 7748
rect 9195 7699 9237 7708
rect 8043 7664 8085 7673
rect 8043 7624 8044 7664
rect 8084 7624 8085 7664
rect 8043 7615 8085 7624
rect 8236 7614 8276 7699
rect 8811 7580 8853 7589
rect 8811 7540 8812 7580
rect 8852 7540 8853 7580
rect 8811 7531 8853 7540
rect 7948 7244 7988 7253
rect 7948 6329 7988 7204
rect 8812 7244 8852 7531
rect 9196 7328 9236 7699
rect 9196 7279 9236 7288
rect 8812 7195 8852 7204
rect 8331 6488 8373 6497
rect 8331 6448 8332 6488
rect 8372 6448 8373 6488
rect 8331 6439 8373 6448
rect 8811 6488 8853 6497
rect 8811 6448 8812 6488
rect 8852 6448 8853 6488
rect 8811 6439 8853 6448
rect 8044 6404 8084 6413
rect 7947 6320 7989 6329
rect 7947 6280 7948 6320
rect 7988 6280 7989 6320
rect 7947 6271 7989 6280
rect 8044 6245 8084 6364
rect 8140 6404 8180 6413
rect 8043 6236 8085 6245
rect 8043 6196 8044 6236
rect 8084 6196 8085 6236
rect 8043 6187 8085 6196
rect 8140 5909 8180 6364
rect 8332 6354 8372 6439
rect 8523 6320 8565 6329
rect 8523 6280 8524 6320
rect 8564 6280 8565 6320
rect 8523 6271 8565 6280
rect 8139 5900 8181 5909
rect 8139 5860 8140 5900
rect 8180 5860 8181 5900
rect 8139 5851 8181 5860
rect 7947 5732 7989 5741
rect 7947 5692 7948 5732
rect 7988 5692 7989 5732
rect 7947 5683 7989 5692
rect 8140 5732 8180 5743
rect 7851 5648 7893 5657
rect 7851 5608 7852 5648
rect 7892 5608 7893 5648
rect 7851 5599 7893 5608
rect 7948 5598 7988 5683
rect 8140 5657 8180 5692
rect 8235 5732 8277 5741
rect 8428 5732 8468 5741
rect 8235 5692 8236 5732
rect 8276 5692 8277 5732
rect 8235 5683 8277 5692
rect 8332 5692 8428 5732
rect 8139 5648 8181 5657
rect 8139 5608 8140 5648
rect 8180 5608 8181 5648
rect 8139 5599 8181 5608
rect 8236 5598 8276 5683
rect 7467 5564 7509 5573
rect 7467 5524 7468 5564
rect 7508 5524 7509 5564
rect 7467 5515 7509 5524
rect 8332 5228 8372 5692
rect 8428 5683 8468 5692
rect 8427 5480 8469 5489
rect 8427 5440 8428 5480
rect 8468 5440 8469 5480
rect 8427 5431 8469 5440
rect 8428 5346 8468 5431
rect 8332 5188 8468 5228
rect 8331 5060 8373 5069
rect 8331 5020 8332 5060
rect 8372 5020 8373 5060
rect 8331 5011 8373 5020
rect 8332 4926 8372 5011
rect 7852 4892 7892 4901
rect 7467 4724 7509 4733
rect 7467 4684 7468 4724
rect 7508 4684 7509 4724
rect 7467 4675 7509 4684
rect 7371 4304 7413 4313
rect 7371 4264 7372 4304
rect 7412 4264 7413 4304
rect 7371 4255 7413 4264
rect 7124 4180 7316 4220
rect 7468 4220 7508 4675
rect 7852 4397 7892 4852
rect 8043 4892 8085 4901
rect 8043 4852 8044 4892
rect 8084 4852 8085 4892
rect 8043 4843 8085 4852
rect 7851 4388 7893 4397
rect 7851 4348 7852 4388
rect 7892 4348 7893 4388
rect 7851 4339 7893 4348
rect 7084 4171 7124 4180
rect 7468 4171 7508 4180
rect 6699 4052 6741 4061
rect 6699 4012 6700 4052
rect 6740 4012 6741 4052
rect 6699 4003 6741 4012
rect 6219 3800 6261 3809
rect 6219 3760 6220 3800
rect 6260 3760 6261 3800
rect 6219 3751 6261 3760
rect 6123 3716 6165 3725
rect 6123 3676 6124 3716
rect 6164 3676 6165 3716
rect 6123 3667 6165 3676
rect 5876 3340 6068 3380
rect 6700 3380 6740 4003
rect 7851 3800 7893 3809
rect 7851 3760 7852 3800
rect 7892 3760 7893 3800
rect 7851 3751 7893 3760
rect 7852 3632 7892 3751
rect 7852 3583 7892 3592
rect 8044 3632 8084 4843
rect 8428 4397 8468 5188
rect 8427 4388 8469 4397
rect 8427 4348 8428 4388
rect 8468 4348 8469 4388
rect 8427 4339 8469 4348
rect 8332 4220 8372 4229
rect 8524 4220 8564 6271
rect 8812 5816 8852 6439
rect 9484 6404 9524 8119
rect 10156 7916 10196 7925
rect 9963 7664 10005 7673
rect 9963 7624 9964 7664
rect 10004 7624 10005 7664
rect 9963 7615 10005 7624
rect 9964 7412 10004 7615
rect 9964 7363 10004 7372
rect 10059 7244 10101 7253
rect 10059 7204 10060 7244
rect 10100 7204 10101 7244
rect 10059 7195 10101 7204
rect 10060 7110 10100 7195
rect 10156 6572 10196 7876
rect 10444 7244 10484 7253
rect 10540 7244 10580 8548
rect 11115 8000 11157 8009
rect 11115 7960 11116 8000
rect 11156 7960 11157 8000
rect 11115 7951 11157 7960
rect 10923 7496 10965 7505
rect 10923 7456 10924 7496
rect 10964 7456 10965 7496
rect 10923 7447 10965 7456
rect 10484 7204 10580 7244
rect 10635 7244 10677 7253
rect 10635 7204 10636 7244
rect 10676 7204 10677 7244
rect 10444 7195 10484 7204
rect 10635 7195 10677 7204
rect 10636 7110 10676 7195
rect 10924 6656 10964 7447
rect 10924 6607 10964 6616
rect 11116 6656 11156 7951
rect 11212 7244 11252 8716
rect 11308 8168 11348 10228
rect 11403 8840 11445 8849
rect 11403 8800 11404 8840
rect 11444 8800 11445 8840
rect 11403 8791 11445 8800
rect 11308 8119 11348 8128
rect 11308 7244 11348 7253
rect 11212 7204 11308 7244
rect 11308 7195 11348 7204
rect 11116 6607 11156 6616
rect 9484 6355 9524 6364
rect 10060 6532 10156 6572
rect 10060 6329 10100 6532
rect 10156 6523 10196 6532
rect 10732 6488 10772 6497
rect 11308 6488 11348 6497
rect 11404 6488 11444 8791
rect 10772 6448 11252 6488
rect 10732 6439 10772 6448
rect 10059 6320 10101 6329
rect 10059 6280 10060 6320
rect 10100 6280 10101 6320
rect 10059 6271 10101 6280
rect 11115 6320 11157 6329
rect 11115 6280 11116 6320
rect 11156 6280 11157 6320
rect 11115 6271 11157 6280
rect 8812 5767 8852 5776
rect 8620 5732 8660 5741
rect 8620 5069 8660 5692
rect 9195 5732 9237 5741
rect 9195 5692 9196 5732
rect 9236 5692 9237 5732
rect 9195 5683 9237 5692
rect 10060 5732 10100 6271
rect 10060 5683 10100 5692
rect 9196 5598 9236 5683
rect 8619 5060 8661 5069
rect 8619 5020 8620 5060
rect 8660 5020 8661 5060
rect 8619 5011 8661 5020
rect 11116 5060 11156 6271
rect 11212 5900 11252 6448
rect 11348 6448 11444 6488
rect 11308 6439 11348 6448
rect 11307 6320 11349 6329
rect 11307 6280 11308 6320
rect 11348 6280 11349 6320
rect 11307 6271 11349 6280
rect 11212 5851 11252 5860
rect 11116 5011 11156 5020
rect 11308 4976 11348 6271
rect 11308 4927 11348 4936
rect 9004 4892 9044 4901
rect 9044 4852 9524 4892
rect 9004 4843 9044 4852
rect 8715 4388 8757 4397
rect 8715 4348 8716 4388
rect 8756 4348 8757 4388
rect 8715 4339 8757 4348
rect 9484 4388 9524 4852
rect 9484 4339 9524 4348
rect 8372 4180 8564 4220
rect 8332 4171 8372 4180
rect 8716 3809 8756 4339
rect 8715 3800 8757 3809
rect 8715 3760 8716 3800
rect 8756 3760 8757 3800
rect 8715 3751 8757 3760
rect 8044 3583 8084 3592
rect 5452 3331 5492 3340
rect 5836 3331 5876 3340
rect 6700 3331 6740 3340
rect 8716 3380 8756 3751
rect 8908 3548 8948 3557
rect 8908 3389 8948 3508
rect 9100 3464 9140 3473
rect 8716 3331 8756 3340
rect 8907 3380 8949 3389
rect 8907 3340 8908 3380
rect 8948 3340 8949 3380
rect 8907 3331 8949 3340
rect 5260 3246 5300 3331
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 9100 1289 9140 3424
rect 6987 1280 7029 1289
rect 6987 1240 6988 1280
rect 7028 1240 7029 1280
rect 6987 1231 7029 1240
rect 9099 1280 9141 1289
rect 9099 1240 9100 1280
rect 9140 1240 9141 1280
rect 9099 1231 9141 1240
rect 6988 80 7028 1231
rect 6968 0 7048 80
<< via2 >>
rect 2860 13840 2900 13880
rect 4108 13840 4148 13880
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 3148 12580 3188 12620
rect 5068 12580 5108 12620
rect 5932 12580 5972 12620
rect 1900 11908 1940 11948
rect 3052 11908 3092 11948
rect 2380 11740 2420 11780
rect 2860 11740 2900 11780
rect 3340 12496 3380 12536
rect 3628 12496 3668 12536
rect 4588 12496 4628 12536
rect 4876 12496 4916 12536
rect 3244 12412 3284 12452
rect 4396 12328 4436 12368
rect 3820 12244 3860 12284
rect 4300 11908 4340 11948
rect 3532 11824 3572 11864
rect 4012 11824 4052 11864
rect 3436 11740 3476 11780
rect 1708 11488 1748 11528
rect 1228 11320 1268 11360
rect 1420 11320 1460 11360
rect 1228 9136 1268 9176
rect 1516 8800 1556 8840
rect 1420 8716 1460 8756
rect 2188 8800 2228 8840
rect 2956 11656 2996 11696
rect 2956 11320 2996 11360
rect 2764 10060 2804 10100
rect 3916 11656 3956 11696
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 3340 10144 3380 10184
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 4012 9640 4052 9680
rect 3052 9472 3092 9512
rect 1324 8632 1364 8672
rect 1708 8632 1748 8672
rect 2380 8632 2420 8672
rect 1228 7540 1268 7580
rect 2860 8800 2900 8840
rect 2764 8716 2804 8756
rect 3148 9388 3188 9428
rect 5356 12412 5396 12452
rect 4972 12328 5012 12368
rect 5452 12244 5492 12284
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 4780 11740 4820 11780
rect 6316 12412 6356 12452
rect 4780 10564 4820 10604
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 5068 10396 5108 10436
rect 4396 10228 4436 10268
rect 5356 10228 5396 10268
rect 5260 10060 5300 10100
rect 4492 9472 4532 9512
rect 4684 9388 4724 9428
rect 5644 9556 5684 9596
rect 3244 8800 3284 8840
rect 3340 8632 3380 8672
rect 1420 7708 1460 7748
rect 1900 7708 1940 7748
rect 1132 6952 1172 6992
rect 1228 6364 1268 6404
rect 1612 7120 1652 7160
rect 1996 7288 2036 7328
rect 1708 7036 1748 7076
rect 2092 7036 2132 7076
rect 1420 5944 1460 5984
rect 1612 5776 1652 5816
rect 1324 5692 1364 5732
rect 2284 6364 2324 6404
rect 2476 6364 2516 6404
rect 2092 5692 2132 5732
rect 2572 5692 2612 5732
rect 3436 7540 3476 7580
rect 2860 5776 2900 5816
rect 3340 7204 3380 7244
rect 3244 7036 3284 7076
rect 4108 8716 4148 8756
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4492 8884 4532 8924
rect 4492 8716 4532 8756
rect 4300 8548 4340 8588
rect 4204 7876 4244 7916
rect 4300 7624 4340 7664
rect 3820 7372 3860 7412
rect 3820 7204 3860 7244
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 2956 5608 2996 5648
rect 3148 5692 3188 5732
rect 4396 7540 4436 7580
rect 4588 8632 4628 8672
rect 4588 7876 4628 7916
rect 4492 7204 4532 7244
rect 4396 6952 4436 6992
rect 4300 5944 4340 5984
rect 3820 5860 3860 5900
rect 4684 7708 4724 7748
rect 4684 7372 4724 7412
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 5068 8884 5108 8924
rect 4972 8296 5012 8336
rect 5452 8548 5492 8588
rect 5260 7792 5300 7832
rect 4876 7708 4916 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 5356 7540 5396 7580
rect 5068 7372 5108 7412
rect 4972 7204 5012 7244
rect 4780 6364 4820 6404
rect 5644 8296 5684 8336
rect 6124 10228 6164 10268
rect 5932 9556 5972 9596
rect 5932 8800 5972 8840
rect 6892 10228 6932 10268
rect 6700 10060 6740 10100
rect 6412 9388 6452 9428
rect 7084 10144 7124 10184
rect 8236 11740 8276 11780
rect 9580 11740 9620 11780
rect 7564 11656 7604 11696
rect 9772 11656 9812 11696
rect 10636 11656 10676 11696
rect 11116 11656 11156 11696
rect 8524 11488 8564 11528
rect 9964 11488 10004 11528
rect 7660 10396 7700 10436
rect 8044 10396 8084 10436
rect 7660 10144 7700 10184
rect 7372 10060 7412 10100
rect 7660 9892 7700 9932
rect 6988 9472 7028 9512
rect 6796 9388 6836 9428
rect 6604 8632 6644 8672
rect 6124 8548 6164 8588
rect 6412 7876 6452 7916
rect 5836 7792 5876 7832
rect 8140 9892 8180 9932
rect 7948 9388 7988 9428
rect 7948 9220 7988 9260
rect 8620 9388 8660 9428
rect 9004 9220 9044 9260
rect 7468 8800 7508 8840
rect 7852 8800 7892 8840
rect 6988 8548 7028 8588
rect 7564 8548 7604 8588
rect 7084 8128 7124 8168
rect 5932 6364 5972 6404
rect 4684 5860 4724 5900
rect 3532 5692 3572 5732
rect 4588 5692 4628 5732
rect 5644 6280 5684 6320
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 4876 5692 4916 5732
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 3340 5020 3380 5060
rect 3148 4936 3188 4976
rect 3052 4852 3092 4892
rect 3436 4852 3476 4892
rect 4300 4852 4340 4892
rect 4588 4852 4628 4892
rect 4588 4096 4628 4136
rect 5452 5440 5492 5480
rect 5260 5020 5300 5060
rect 4780 4852 4820 4892
rect 5068 4684 5108 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 5356 4516 5396 4556
rect 5068 4348 5108 4388
rect 4780 4264 4820 4304
rect 5260 4264 5300 4304
rect 5548 4684 5588 4724
rect 5164 4096 5204 4136
rect 3916 4012 3956 4052
rect 4684 4012 4724 4052
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 3244 3676 3284 3716
rect 5068 3424 5108 3464
rect 5260 3340 5300 3380
rect 6892 5860 6932 5900
rect 6604 5692 6644 5732
rect 5932 5608 5972 5648
rect 6220 5608 6260 5648
rect 5932 4768 5972 4808
rect 5644 3424 5684 3464
rect 6412 5440 6452 5480
rect 6412 5020 6452 5060
rect 6220 4684 6260 4724
rect 6316 4348 6356 4388
rect 6796 5440 6836 5480
rect 6700 4852 6740 4892
rect 6700 4432 6740 4472
rect 8908 8800 8948 8840
rect 8428 8548 8468 8588
rect 7564 6364 7604 6404
rect 7372 6280 7412 6320
rect 7468 6196 7508 6236
rect 7084 5776 7124 5816
rect 7084 5524 7124 5564
rect 7180 4432 7220 4472
rect 7948 7960 7988 8000
rect 8332 7876 8372 7916
rect 9100 8716 9140 8756
rect 9004 8632 9044 8672
rect 8908 8464 8948 8504
rect 8524 7960 8564 8000
rect 8716 7960 8756 8000
rect 10444 10228 10484 10268
rect 9388 10060 9428 10100
rect 11020 10228 11060 10268
rect 9964 8716 10004 8756
rect 10156 8632 10196 8672
rect 11116 8800 11156 8840
rect 9292 8464 9332 8504
rect 9196 8128 9236 8168
rect 9484 8128 9524 8168
rect 9292 7876 9332 7916
rect 8236 7708 8276 7748
rect 9196 7708 9236 7748
rect 8044 7624 8084 7664
rect 8812 7540 8852 7580
rect 8332 6448 8372 6488
rect 8812 6448 8852 6488
rect 7948 6280 7988 6320
rect 8044 6196 8084 6236
rect 8524 6280 8564 6320
rect 8140 5860 8180 5900
rect 7948 5692 7988 5732
rect 7852 5608 7892 5648
rect 8236 5692 8276 5732
rect 8140 5608 8180 5648
rect 7468 5524 7508 5564
rect 8428 5440 8468 5480
rect 8332 5020 8372 5060
rect 7468 4684 7508 4724
rect 7372 4264 7412 4304
rect 8044 4852 8084 4892
rect 7852 4348 7892 4388
rect 6700 4012 6740 4052
rect 6220 3760 6260 3800
rect 6124 3676 6164 3716
rect 7852 3760 7892 3800
rect 8428 4348 8468 4388
rect 9964 7624 10004 7664
rect 10060 7204 10100 7244
rect 11116 7960 11156 8000
rect 10924 7456 10964 7496
rect 10636 7204 10676 7244
rect 11404 8800 11444 8840
rect 10060 6280 10100 6320
rect 11116 6280 11156 6320
rect 9196 5692 9236 5732
rect 8620 5020 8660 5060
rect 11308 6280 11348 6320
rect 8716 4348 8756 4388
rect 8716 3760 8756 3800
rect 8908 3340 8948 3380
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 6988 1240 7028 1280
rect 9100 1240 9140 1280
<< metal3 >>
rect 2851 13840 2860 13880
rect 2900 13840 4108 13880
rect 4148 13840 4157 13880
rect 3679 12832 3688 12872
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 4056 12832 4065 12872
rect 3139 12580 3148 12620
rect 3188 12580 5068 12620
rect 5108 12580 5932 12620
rect 5972 12580 5981 12620
rect 3331 12496 3340 12536
rect 3380 12496 3628 12536
rect 3668 12496 4588 12536
rect 4628 12496 4876 12536
rect 4916 12496 4925 12536
rect 6307 12452 6365 12453
rect 3235 12412 3244 12452
rect 3284 12412 5356 12452
rect 5396 12412 5405 12452
rect 6222 12412 6316 12452
rect 6356 12412 6365 12452
rect 6307 12411 6365 12412
rect 4387 12328 4396 12368
rect 4436 12328 4972 12368
rect 5012 12328 5021 12368
rect 3811 12244 3820 12284
rect 3860 12244 5452 12284
rect 5492 12244 5501 12284
rect 4919 12076 4928 12116
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 5296 12076 5305 12116
rect 1891 11948 1949 11949
rect 1806 11908 1900 11948
rect 1940 11908 1949 11948
rect 3043 11908 3052 11948
rect 3092 11908 4300 11948
rect 4340 11908 4349 11948
rect 1891 11907 1949 11908
rect 3523 11824 3532 11864
rect 3572 11824 4012 11864
rect 4052 11824 4061 11864
rect 2371 11740 2380 11780
rect 2420 11740 2860 11780
rect 2900 11740 2909 11780
rect 3427 11740 3436 11780
rect 3476 11740 4780 11780
rect 4820 11740 4829 11780
rect 8227 11740 8236 11780
rect 8276 11740 9580 11780
rect 9620 11740 9629 11780
rect 2947 11656 2956 11696
rect 2996 11656 3916 11696
rect 3956 11656 3965 11696
rect 7555 11656 7564 11696
rect 7604 11656 9772 11696
rect 9812 11656 10636 11696
rect 10676 11656 11116 11696
rect 11156 11656 11165 11696
rect 0 11528 80 11548
rect 0 11488 1708 11528
rect 1748 11488 1757 11528
rect 8515 11488 8524 11528
rect 8564 11488 9964 11528
rect 10004 11488 10013 11528
rect 0 11468 80 11488
rect 2500 11404 2996 11444
rect 0 11360 80 11380
rect 0 11320 500 11360
rect 1219 11320 1228 11360
rect 1268 11320 1277 11360
rect 1411 11320 1420 11360
rect 1460 11320 1469 11360
rect 0 11300 80 11320
rect 460 11276 500 11320
rect 1228 11276 1268 11320
rect 460 11236 1268 11276
rect 1420 11276 1460 11320
rect 2500 11276 2540 11404
rect 2956 11360 2996 11404
rect 2916 11320 2956 11360
rect 2996 11320 3005 11360
rect 3679 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 4065 11360
rect 1420 11236 2540 11276
rect 4771 10564 4780 10604
rect 4820 10564 4829 10604
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 4780 10436 4820 10564
rect 4780 10396 5068 10436
rect 5108 10396 5117 10436
rect 7651 10396 7660 10436
rect 7700 10396 8044 10436
rect 8084 10396 8093 10436
rect 4387 10228 4396 10268
rect 4436 10228 5356 10268
rect 5396 10228 5405 10268
rect 6115 10228 6124 10268
rect 6164 10228 6892 10268
rect 6932 10228 6941 10268
rect 10435 10228 10444 10268
rect 10484 10228 11020 10268
rect 11060 10228 11069 10268
rect 3331 10144 3340 10184
rect 3380 10144 5300 10184
rect 7075 10144 7084 10184
rect 7124 10144 7660 10184
rect 7700 10144 7709 10184
rect 5260 10100 5300 10144
rect 2755 10060 2764 10100
rect 2804 10060 4148 10100
rect 5251 10060 5260 10100
rect 5300 10060 5309 10100
rect 6691 10060 6700 10100
rect 6740 10060 7372 10100
rect 7412 10060 9388 10100
rect 9428 10060 9437 10100
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 4108 9680 4148 10060
rect 7651 9892 7660 9932
rect 7700 9892 8140 9932
rect 8180 9892 8189 9932
rect 4003 9640 4012 9680
rect 4052 9640 4148 9680
rect 5635 9556 5644 9596
rect 5684 9556 5932 9596
rect 5972 9556 5981 9596
rect 3043 9472 3052 9512
rect 3092 9472 4492 9512
rect 4532 9472 6988 9512
rect 7028 9472 7037 9512
rect 3139 9388 3148 9428
rect 3188 9388 4684 9428
rect 4724 9388 6412 9428
rect 6452 9388 6796 9428
rect 6836 9388 6845 9428
rect 7939 9388 7948 9428
rect 7988 9388 8620 9428
rect 8660 9388 8669 9428
rect 7939 9220 7948 9260
rect 7988 9220 9004 9260
rect 9044 9220 9053 9260
rect 0 9176 80 9196
rect 0 9136 1228 9176
rect 1268 9136 1277 9176
rect 0 9116 80 9136
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 4483 8884 4492 8924
rect 4532 8884 5068 8924
rect 5108 8884 5117 8924
rect 12504 8840 12584 8860
rect 1507 8800 1516 8840
rect 1556 8800 2188 8840
rect 2228 8800 2860 8840
rect 2900 8800 2909 8840
rect 3235 8800 3244 8840
rect 3284 8800 5932 8840
rect 5972 8800 5981 8840
rect 7459 8800 7468 8840
rect 7508 8800 7852 8840
rect 7892 8800 7901 8840
rect 8899 8800 8908 8840
rect 8948 8800 11116 8840
rect 11156 8800 11165 8840
rect 11395 8800 11404 8840
rect 11444 8800 12584 8840
rect 12504 8780 12584 8800
rect 1411 8716 1420 8756
rect 1460 8716 2764 8756
rect 2804 8716 2813 8756
rect 4099 8716 4108 8756
rect 4148 8716 4492 8756
rect 4532 8716 4541 8756
rect 9091 8716 9100 8756
rect 9140 8716 9964 8756
rect 10004 8716 10013 8756
rect 1315 8632 1324 8672
rect 1364 8632 1708 8672
rect 1748 8632 2380 8672
rect 2420 8632 2540 8672
rect 3331 8632 3340 8672
rect 3380 8632 4588 8672
rect 4628 8632 6604 8672
rect 6644 8632 6653 8672
rect 8995 8632 9004 8672
rect 9044 8632 10156 8672
rect 10196 8632 10205 8672
rect 2500 8588 2540 8632
rect 2500 8548 4300 8588
rect 4340 8548 5452 8588
rect 5492 8548 6124 8588
rect 6164 8548 6173 8588
rect 6979 8548 6988 8588
rect 7028 8548 7564 8588
rect 7604 8548 8428 8588
rect 8468 8548 8477 8588
rect 8899 8464 8908 8504
rect 8948 8464 9292 8504
rect 9332 8464 9341 8504
rect 5347 8336 5405 8337
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 4963 8296 4972 8336
rect 5012 8296 5356 8336
rect 5396 8296 5644 8336
rect 5684 8296 5693 8336
rect 5347 8295 5405 8296
rect 7075 8128 7084 8168
rect 7124 8128 9196 8168
rect 9236 8128 9484 8168
rect 9524 8128 9533 8168
rect 7939 7960 7948 8000
rect 7988 7960 8524 8000
rect 8564 7960 8573 8000
rect 8707 7960 8716 8000
rect 8756 7960 11116 8000
rect 11156 7960 11165 8000
rect 4195 7876 4204 7916
rect 4244 7876 4588 7916
rect 4628 7876 6412 7916
rect 6452 7876 6461 7916
rect 8323 7876 8332 7916
rect 8372 7876 9292 7916
rect 9332 7876 9341 7916
rect 5251 7792 5260 7832
rect 5300 7792 5836 7832
rect 5876 7792 5885 7832
rect 1411 7708 1420 7748
rect 1460 7708 1900 7748
rect 1940 7708 4684 7748
rect 4724 7708 4733 7748
rect 4867 7708 4876 7748
rect 4916 7708 4925 7748
rect 8227 7708 8236 7748
rect 8276 7708 9196 7748
rect 9236 7708 9245 7748
rect 4876 7664 4916 7708
rect 4291 7624 4300 7664
rect 4340 7624 4916 7664
rect 8035 7624 8044 7664
rect 8084 7624 9964 7664
rect 10004 7624 10013 7664
rect 1219 7540 1228 7580
rect 1268 7540 3436 7580
rect 3476 7540 3485 7580
rect 4387 7540 4396 7580
rect 4436 7540 4820 7580
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 5347 7540 5356 7580
rect 5396 7540 8812 7580
rect 8852 7540 8861 7580
rect 4780 7412 4820 7540
rect 12504 7496 12584 7516
rect 10915 7456 10924 7496
rect 10964 7456 12584 7496
rect 12504 7436 12584 7456
rect 3811 7372 3820 7412
rect 3860 7372 4684 7412
rect 4724 7372 4733 7412
rect 4780 7372 5068 7412
rect 5108 7372 5117 7412
rect 1987 7288 1996 7328
rect 2036 7288 4532 7328
rect 4492 7244 4532 7288
rect 5347 7244 5405 7245
rect 3331 7204 3340 7244
rect 3380 7204 3820 7244
rect 3860 7204 3869 7244
rect 4483 7204 4492 7244
rect 4532 7204 4541 7244
rect 4963 7204 4972 7244
rect 5012 7204 5356 7244
rect 5396 7204 5405 7244
rect 10051 7204 10060 7244
rect 10100 7204 10636 7244
rect 10676 7204 10685 7244
rect 5347 7203 5405 7204
rect 1603 7120 1612 7160
rect 1652 7120 3284 7160
rect 3244 7076 3284 7120
rect 1699 7036 1708 7076
rect 1748 7036 2092 7076
rect 2132 7036 2540 7076
rect 3235 7036 3244 7076
rect 3284 7036 3293 7076
rect 0 6992 80 7012
rect 2500 6992 2540 7036
rect 0 6952 1132 6992
rect 1172 6952 1181 6992
rect 2500 6952 4396 6992
rect 4436 6952 4445 6992
rect 0 6932 80 6952
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 8323 6448 8332 6488
rect 8372 6448 8812 6488
rect 8852 6448 8861 6488
rect 1219 6364 1228 6404
rect 1268 6364 2284 6404
rect 2324 6364 2333 6404
rect 2467 6364 2476 6404
rect 2516 6364 4780 6404
rect 4820 6364 5932 6404
rect 5972 6364 5981 6404
rect 7555 6364 7564 6404
rect 7604 6364 11156 6404
rect 11116 6320 11156 6364
rect 12504 6320 12584 6340
rect 5635 6280 5644 6320
rect 5684 6280 7372 6320
rect 7412 6280 7421 6320
rect 7939 6280 7948 6320
rect 7988 6280 8524 6320
rect 8564 6280 10060 6320
rect 10100 6280 10109 6320
rect 11107 6280 11116 6320
rect 11156 6280 11165 6320
rect 11299 6280 11308 6320
rect 11348 6280 12584 6320
rect 12504 6260 12584 6280
rect 7459 6196 7468 6236
rect 7508 6196 8044 6236
rect 8084 6196 8093 6236
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 1411 5944 1420 5984
rect 1460 5944 4300 5984
rect 4340 5944 4349 5984
rect 3811 5860 3820 5900
rect 3860 5860 4684 5900
rect 4724 5860 4733 5900
rect 6883 5860 6892 5900
rect 6932 5860 8140 5900
rect 8180 5860 8189 5900
rect 0 5816 80 5836
rect 0 5776 1612 5816
rect 1652 5776 1661 5816
rect 2851 5776 2860 5816
rect 2900 5776 7084 5816
rect 7124 5776 7133 5816
rect 0 5756 80 5776
rect 1315 5692 1324 5732
rect 1364 5692 2092 5732
rect 2132 5692 2141 5732
rect 2563 5692 2572 5732
rect 2612 5692 3148 5732
rect 3188 5692 3532 5732
rect 3572 5692 3581 5732
rect 4579 5692 4588 5732
rect 4628 5692 4876 5732
rect 4916 5692 4925 5732
rect 6595 5692 6604 5732
rect 6644 5692 7948 5732
rect 7988 5692 7997 5732
rect 8227 5692 8236 5732
rect 8276 5692 9196 5732
rect 9236 5692 9245 5732
rect 2947 5608 2956 5648
rect 2996 5608 5932 5648
rect 5972 5608 5981 5648
rect 6211 5608 6220 5648
rect 6260 5608 7852 5648
rect 7892 5608 8140 5648
rect 8180 5608 8189 5648
rect 7075 5524 7084 5564
rect 7124 5524 7468 5564
rect 7508 5524 7517 5564
rect 5443 5440 5452 5480
rect 5492 5440 6412 5480
rect 6452 5440 6461 5480
rect 6787 5440 6796 5480
rect 6836 5440 8428 5480
rect 8468 5440 8477 5480
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 3331 5020 3340 5060
rect 3380 5020 5260 5060
rect 5300 5020 5309 5060
rect 6403 5020 6412 5060
rect 6452 5020 8332 5060
rect 8372 5020 8620 5060
rect 8660 5020 8669 5060
rect 3139 4936 3148 4976
rect 3188 4936 4628 4976
rect 4588 4892 4628 4936
rect 3043 4852 3052 4892
rect 3092 4852 3101 4892
rect 3427 4852 3436 4892
rect 3476 4852 4300 4892
rect 4340 4852 4349 4892
rect 4579 4852 4588 4892
rect 4628 4852 4780 4892
rect 4820 4852 4829 4892
rect 6691 4852 6700 4892
rect 6740 4852 8044 4892
rect 8084 4852 8093 4892
rect 3052 4808 3092 4852
rect 3052 4768 5932 4808
rect 5972 4768 5981 4808
rect 5059 4684 5068 4724
rect 5108 4684 5548 4724
rect 5588 4684 5597 4724
rect 6211 4684 6220 4724
rect 6260 4684 7468 4724
rect 7508 4684 7517 4724
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 5347 4516 5356 4556
rect 5396 4516 5405 4556
rect 5356 4388 5396 4516
rect 6691 4432 6700 4472
rect 6740 4432 7180 4472
rect 7220 4432 7229 4472
rect 5059 4348 5068 4388
rect 5108 4348 5396 4388
rect 6307 4348 6316 4388
rect 6356 4348 7852 4388
rect 7892 4348 7901 4388
rect 8419 4348 8428 4388
rect 8468 4348 8716 4388
rect 8756 4348 8765 4388
rect 12504 4304 12584 4324
rect 4771 4264 4780 4304
rect 4820 4264 5260 4304
rect 5300 4264 5309 4304
rect 7363 4264 7372 4304
rect 7412 4264 12584 4304
rect 12504 4244 12584 4264
rect 4579 4096 4588 4136
rect 4628 4096 5164 4136
rect 5204 4096 5213 4136
rect 3907 4012 3916 4052
rect 3956 4012 4684 4052
rect 4724 4012 6700 4052
rect 6740 4012 6749 4052
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 6211 3760 6220 3800
rect 6260 3760 7852 3800
rect 7892 3760 8716 3800
rect 8756 3760 8765 3800
rect 3235 3676 3244 3716
rect 3284 3676 6124 3716
rect 6164 3676 6173 3716
rect 5059 3424 5068 3464
rect 5108 3424 5644 3464
rect 5684 3424 5693 3464
rect 5251 3340 5260 3380
rect 5300 3340 8908 3380
rect 8948 3340 8957 3380
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 6979 1240 6988 1280
rect 7028 1240 9100 1280
rect 9140 1240 9149 1280
<< via3 >>
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 6316 12412 6356 12452
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 1900 11908 1940 11948
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 5356 8296 5396 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 5356 7204 5396 7244
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
<< metal4 >>
rect 3688 12872 4056 12881
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 3688 12823 4056 12832
rect 1899 12452 1941 12461
rect 1899 12412 1900 12452
rect 1940 12412 1941 12452
rect 1899 12403 1941 12412
rect 6315 12452 6357 12461
rect 6315 12412 6316 12452
rect 6356 12412 6357 12452
rect 6315 12403 6357 12412
rect 1900 11948 1940 12403
rect 6316 12318 6356 12403
rect 4928 12116 5296 12125
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 4928 12067 5296 12076
rect 1900 11899 1940 11908
rect 3688 11360 4056 11369
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 3688 11311 4056 11320
rect 4928 10604 5296 10613
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 4928 10555 5296 10564
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 5356 8336 5396 8345
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 5356 7244 5396 8296
rect 5356 7195 5396 7204
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
<< via4 >>
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 1900 12412 1940 12452
rect 6316 12412 6356 12452
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
<< metal5 >>
rect 3679 12872 3726 12914
rect 3850 12872 3894 12914
rect 4018 12872 4065 12914
rect 3679 12832 3688 12872
rect 3850 12832 3852 12872
rect 3892 12832 3894 12872
rect 4056 12832 4065 12872
rect 3679 12790 3726 12832
rect 3850 12790 3894 12832
rect 4018 12790 4065 12832
rect 1891 12412 1900 12452
rect 1940 12412 6316 12452
rect 6356 12412 6365 12452
rect 4919 12116 4966 12158
rect 5090 12116 5134 12158
rect 5258 12116 5305 12158
rect 4919 12076 4928 12116
rect 5090 12076 5092 12116
rect 5132 12076 5134 12116
rect 5296 12076 5305 12116
rect 4919 12034 4966 12076
rect 5090 12034 5134 12076
rect 5258 12034 5305 12076
rect 3679 11360 3726 11402
rect 3850 11360 3894 11402
rect 4018 11360 4065 11402
rect 3679 11320 3688 11360
rect 3850 11320 3852 11360
rect 3892 11320 3894 11360
rect 4056 11320 4065 11360
rect 3679 11278 3726 11320
rect 3850 11278 3894 11320
rect 4018 11278 4065 11320
rect 4919 10604 4966 10646
rect 5090 10604 5134 10646
rect 5258 10604 5305 10646
rect 4919 10564 4928 10604
rect 5090 10564 5092 10604
rect 5132 10564 5134 10604
rect 5296 10564 5305 10604
rect 4919 10522 4966 10564
rect 5090 10522 5134 10564
rect 5258 10522 5305 10564
rect 3679 9848 3726 9890
rect 3850 9848 3894 9890
rect 4018 9848 4065 9890
rect 3679 9808 3688 9848
rect 3850 9808 3852 9848
rect 3892 9808 3894 9848
rect 4056 9808 4065 9848
rect 3679 9766 3726 9808
rect 3850 9766 3894 9808
rect 4018 9766 4065 9808
rect 4919 9092 4966 9134
rect 5090 9092 5134 9134
rect 5258 9092 5305 9134
rect 4919 9052 4928 9092
rect 5090 9052 5092 9092
rect 5132 9052 5134 9092
rect 5296 9052 5305 9092
rect 4919 9010 4966 9052
rect 5090 9010 5134 9052
rect 5258 9010 5305 9052
rect 3679 8336 3726 8378
rect 3850 8336 3894 8378
rect 4018 8336 4065 8378
rect 3679 8296 3688 8336
rect 3850 8296 3852 8336
rect 3892 8296 3894 8336
rect 4056 8296 4065 8336
rect 3679 8254 3726 8296
rect 3850 8254 3894 8296
rect 4018 8254 4065 8296
rect 4919 7580 4966 7622
rect 5090 7580 5134 7622
rect 5258 7580 5305 7622
rect 4919 7540 4928 7580
rect 5090 7540 5092 7580
rect 5132 7540 5134 7580
rect 5296 7540 5305 7580
rect 4919 7498 4966 7540
rect 5090 7498 5134 7540
rect 5258 7498 5305 7540
rect 3679 6824 3726 6866
rect 3850 6824 3894 6866
rect 4018 6824 4065 6866
rect 3679 6784 3688 6824
rect 3850 6784 3852 6824
rect 3892 6784 3894 6824
rect 4056 6784 4065 6824
rect 3679 6742 3726 6784
rect 3850 6742 3894 6784
rect 4018 6742 4065 6784
rect 4919 6068 4966 6110
rect 5090 6068 5134 6110
rect 5258 6068 5305 6110
rect 4919 6028 4928 6068
rect 5090 6028 5092 6068
rect 5132 6028 5134 6068
rect 5296 6028 5305 6068
rect 4919 5986 4966 6028
rect 5090 5986 5134 6028
rect 5258 5986 5305 6028
rect 3679 5312 3726 5354
rect 3850 5312 3894 5354
rect 4018 5312 4065 5354
rect 3679 5272 3688 5312
rect 3850 5272 3852 5312
rect 3892 5272 3894 5312
rect 4056 5272 4065 5312
rect 3679 5230 3726 5272
rect 3850 5230 3894 5272
rect 4018 5230 4065 5272
rect 4919 4556 4966 4598
rect 5090 4556 5134 4598
rect 5258 4556 5305 4598
rect 4919 4516 4928 4556
rect 5090 4516 5092 4556
rect 5132 4516 5134 4556
rect 5296 4516 5305 4556
rect 4919 4474 4966 4516
rect 5090 4474 5134 4516
rect 5258 4474 5305 4516
rect 3679 3800 3726 3842
rect 3850 3800 3894 3842
rect 4018 3800 4065 3842
rect 3679 3760 3688 3800
rect 3850 3760 3852 3800
rect 3892 3760 3894 3800
rect 4056 3760 4065 3800
rect 3679 3718 3726 3760
rect 3850 3718 3894 3760
rect 4018 3718 4065 3760
rect 4919 3044 4966 3086
rect 5090 3044 5134 3086
rect 5258 3044 5305 3086
rect 4919 3004 4928 3044
rect 5090 3004 5092 3044
rect 5132 3004 5134 3044
rect 5296 3004 5305 3044
rect 4919 2962 4966 3004
rect 5090 2962 5134 3004
rect 5258 2962 5305 3004
<< via5 >>
rect 3726 12872 3850 12914
rect 3894 12872 4018 12914
rect 3726 12832 3728 12872
rect 3728 12832 3770 12872
rect 3770 12832 3810 12872
rect 3810 12832 3850 12872
rect 3894 12832 3934 12872
rect 3934 12832 3974 12872
rect 3974 12832 4016 12872
rect 4016 12832 4018 12872
rect 3726 12790 3850 12832
rect 3894 12790 4018 12832
rect 4966 12116 5090 12158
rect 5134 12116 5258 12158
rect 4966 12076 4968 12116
rect 4968 12076 5010 12116
rect 5010 12076 5050 12116
rect 5050 12076 5090 12116
rect 5134 12076 5174 12116
rect 5174 12076 5214 12116
rect 5214 12076 5256 12116
rect 5256 12076 5258 12116
rect 4966 12034 5090 12076
rect 5134 12034 5258 12076
rect 3726 11360 3850 11402
rect 3894 11360 4018 11402
rect 3726 11320 3728 11360
rect 3728 11320 3770 11360
rect 3770 11320 3810 11360
rect 3810 11320 3850 11360
rect 3894 11320 3934 11360
rect 3934 11320 3974 11360
rect 3974 11320 4016 11360
rect 4016 11320 4018 11360
rect 3726 11278 3850 11320
rect 3894 11278 4018 11320
rect 4966 10604 5090 10646
rect 5134 10604 5258 10646
rect 4966 10564 4968 10604
rect 4968 10564 5010 10604
rect 5010 10564 5050 10604
rect 5050 10564 5090 10604
rect 5134 10564 5174 10604
rect 5174 10564 5214 10604
rect 5214 10564 5256 10604
rect 5256 10564 5258 10604
rect 4966 10522 5090 10564
rect 5134 10522 5258 10564
rect 3726 9848 3850 9890
rect 3894 9848 4018 9890
rect 3726 9808 3728 9848
rect 3728 9808 3770 9848
rect 3770 9808 3810 9848
rect 3810 9808 3850 9848
rect 3894 9808 3934 9848
rect 3934 9808 3974 9848
rect 3974 9808 4016 9848
rect 4016 9808 4018 9848
rect 3726 9766 3850 9808
rect 3894 9766 4018 9808
rect 4966 9092 5090 9134
rect 5134 9092 5258 9134
rect 4966 9052 4968 9092
rect 4968 9052 5010 9092
rect 5010 9052 5050 9092
rect 5050 9052 5090 9092
rect 5134 9052 5174 9092
rect 5174 9052 5214 9092
rect 5214 9052 5256 9092
rect 5256 9052 5258 9092
rect 4966 9010 5090 9052
rect 5134 9010 5258 9052
rect 3726 8336 3850 8378
rect 3894 8336 4018 8378
rect 3726 8296 3728 8336
rect 3728 8296 3770 8336
rect 3770 8296 3810 8336
rect 3810 8296 3850 8336
rect 3894 8296 3934 8336
rect 3934 8296 3974 8336
rect 3974 8296 4016 8336
rect 4016 8296 4018 8336
rect 3726 8254 3850 8296
rect 3894 8254 4018 8296
rect 4966 7580 5090 7622
rect 5134 7580 5258 7622
rect 4966 7540 4968 7580
rect 4968 7540 5010 7580
rect 5010 7540 5050 7580
rect 5050 7540 5090 7580
rect 5134 7540 5174 7580
rect 5174 7540 5214 7580
rect 5214 7540 5256 7580
rect 5256 7540 5258 7580
rect 4966 7498 5090 7540
rect 5134 7498 5258 7540
rect 3726 6824 3850 6866
rect 3894 6824 4018 6866
rect 3726 6784 3728 6824
rect 3728 6784 3770 6824
rect 3770 6784 3810 6824
rect 3810 6784 3850 6824
rect 3894 6784 3934 6824
rect 3934 6784 3974 6824
rect 3974 6784 4016 6824
rect 4016 6784 4018 6824
rect 3726 6742 3850 6784
rect 3894 6742 4018 6784
rect 4966 6068 5090 6110
rect 5134 6068 5258 6110
rect 4966 6028 4968 6068
rect 4968 6028 5010 6068
rect 5010 6028 5050 6068
rect 5050 6028 5090 6068
rect 5134 6028 5174 6068
rect 5174 6028 5214 6068
rect 5214 6028 5256 6068
rect 5256 6028 5258 6068
rect 4966 5986 5090 6028
rect 5134 5986 5258 6028
rect 3726 5312 3850 5354
rect 3894 5312 4018 5354
rect 3726 5272 3728 5312
rect 3728 5272 3770 5312
rect 3770 5272 3810 5312
rect 3810 5272 3850 5312
rect 3894 5272 3934 5312
rect 3934 5272 3974 5312
rect 3974 5272 4016 5312
rect 4016 5272 4018 5312
rect 3726 5230 3850 5272
rect 3894 5230 4018 5272
rect 4966 4556 5090 4598
rect 5134 4556 5258 4598
rect 4966 4516 4968 4556
rect 4968 4516 5010 4556
rect 5010 4516 5050 4556
rect 5050 4516 5090 4556
rect 5134 4516 5174 4556
rect 5174 4516 5214 4556
rect 5214 4516 5256 4556
rect 5256 4516 5258 4556
rect 4966 4474 5090 4516
rect 5134 4474 5258 4516
rect 3726 3800 3850 3842
rect 3894 3800 4018 3842
rect 3726 3760 3728 3800
rect 3728 3760 3770 3800
rect 3770 3760 3810 3800
rect 3810 3760 3850 3800
rect 3894 3760 3934 3800
rect 3934 3760 3974 3800
rect 3974 3760 4016 3800
rect 4016 3760 4018 3800
rect 3726 3718 3850 3760
rect 3894 3718 4018 3760
rect 4966 3044 5090 3086
rect 5134 3044 5258 3086
rect 4966 3004 4968 3044
rect 4968 3004 5010 3044
rect 5010 3004 5050 3044
rect 5050 3004 5090 3044
rect 5134 3004 5174 3044
rect 5174 3004 5214 3044
rect 5214 3004 5256 3044
rect 5256 3004 5258 3044
rect 4966 2962 5090 3004
rect 5134 2962 5258 3004
<< metal6 >>
rect 3652 12914 4092 12978
rect 3652 12790 3726 12914
rect 3850 12790 3894 12914
rect 4018 12790 4092 12914
rect 3652 11402 4092 12790
rect 3652 11278 3726 11402
rect 3850 11278 3894 11402
rect 4018 11278 4092 11402
rect 3652 9890 4092 11278
rect 3652 9766 3726 9890
rect 3850 9766 3894 9890
rect 4018 9766 4092 9890
rect 3652 8378 4092 9766
rect 3652 8254 3726 8378
rect 3850 8254 3894 8378
rect 4018 8254 4092 8378
rect 3652 6866 4092 8254
rect 3652 6742 3726 6866
rect 3850 6742 3894 6866
rect 4018 6742 4092 6866
rect 3652 5934 4092 6742
rect 3652 5554 3682 5934
rect 4062 5554 4092 5934
rect 3652 5354 4092 5554
rect 3652 5230 3726 5354
rect 3850 5230 3894 5354
rect 4018 5230 4092 5354
rect 3652 3842 4092 5230
rect 3652 3718 3726 3842
rect 3850 3718 3894 3842
rect 4018 3718 4092 3842
rect 3652 2980 4092 3718
rect 4892 12158 5332 12896
rect 4892 12034 4966 12158
rect 5090 12034 5134 12158
rect 5258 12034 5332 12158
rect 4892 10646 5332 12034
rect 4892 10522 4966 10646
rect 5090 10522 5134 10646
rect 5258 10522 5332 10646
rect 4892 9134 5332 10522
rect 4892 9010 4966 9134
rect 5090 9010 5134 9134
rect 5258 9010 5332 9134
rect 4892 7622 5332 9010
rect 4892 7498 4966 7622
rect 5090 7498 5134 7622
rect 5258 7498 5332 7622
rect 4892 7174 5332 7498
rect 4892 6794 4922 7174
rect 5302 6794 5332 7174
rect 4892 6110 5332 6794
rect 4892 5986 4966 6110
rect 5090 5986 5134 6110
rect 5258 5986 5332 6110
rect 4892 4598 5332 5986
rect 4892 4474 4966 4598
rect 5090 4474 5134 4598
rect 5258 4474 5332 4598
rect 4892 3086 5332 4474
rect 4892 2962 4966 3086
rect 5090 2962 5134 3086
rect 5258 2962 5332 3086
rect 4892 2898 5332 2962
<< via6 >>
rect 3682 5554 4062 5934
rect 4922 6794 5302 7174
<< metal7 >>
rect 1108 7174 11468 7204
rect 1108 6794 4922 7174
rect 5302 6794 11468 7174
rect 1108 6764 11468 6794
rect 1108 5934 11468 5964
rect 1108 5554 3682 5934
rect 4062 5554 11468 5934
rect 1108 5524 11468 5554
use sg13g2_inv_1  _054_
timestamp 1676386529
transform 1 0 8064 0 -1 6048
box -48 -56 336 834
use sg13g2_nand2_1  _055_
timestamp 1676560849
transform 1 0 6144 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _056_
timestamp 1676560849
transform -1 0 7680 0 1 6048
box -48 -56 432 834
use sg13g2_nor2_1  _057_
timestamp 1676630787
transform -1 0 8736 0 -1 6048
box -48 -56 432 834
use sg13g2_xor2_1  _058_
timestamp 1677581577
transform 1 0 6336 0 1 4536
box -48 -56 816 834
use sg13g2_o21ai_1  _059_
timestamp 1685182643
transform -1 0 7008 0 -1 4536
box -48 -56 538 834
use sg13g2_xnor2_1  _060_
timestamp 1677520200
transform 1 0 7680 0 1 6048
box -48 -56 816 834
use sg13g2_nand2_1  _061_
timestamp 1676560849
transform 1 0 2688 0 -1 9072
box -48 -56 432 834
use sg13g2_nand2b_1  _062_
timestamp 1676570795
transform -1 0 2400 0 -1 9072
box -48 -56 528 834
use sg13g2_xnor2_1  _063_
timestamp 1677520200
transform -1 0 2016 0 -1 10584
box -48 -56 816 834
use sg13g2_nand2_1  _064_
timestamp 1676560849
transform 1 0 2784 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _065_
timestamp 1676560849
transform -1 0 5376 0 1 3024
box -48 -56 432 834
use sg13g2_nor2_1  _066_
timestamp 1676630787
transform -1 0 3072 0 1 4536
box -48 -56 432 834
use sg13g2_xor2_1  _067_
timestamp 1677581577
transform -1 0 5952 0 -1 4536
box -48 -56 816 834
use sg13g2_o21ai_1  _068_
timestamp 1685182643
transform 1 0 3072 0 1 4536
box -48 -56 538 834
use sg13g2_xnor2_1  _069_
timestamp 1677520200
transform 1 0 4416 0 1 4536
box -48 -56 816 834
use sg13g2_nand2_1  _070_
timestamp 1676560849
transform 1 0 1824 0 -1 7560
box -48 -56 432 834
use sg13g2_nand2_1  _071_
timestamp 1676560849
transform 1 0 2400 0 -1 6048
box -48 -56 432 834
use sg13g2_nor2_1  _072_
timestamp 1676630787
transform -1 0 1824 0 -1 7560
box -48 -56 432 834
use sg13g2_xor2_1  _073_
timestamp 1677581577
transform -1 0 4224 0 -1 9072
box -48 -56 816 834
use sg13g2_o21ai_1  _074_
timestamp 1685182643
transform 1 0 3072 0 -1 7560
box -48 -56 538 834
use sg13g2_xnor2_1  _075_
timestamp 1677520200
transform 1 0 3168 0 -1 6048
box -48 -56 816 834
use sg13g2_nand2_1  _076_
timestamp 1676560849
transform -1 0 6720 0 1 9072
box -48 -56 432 834
use sg13g2_nand2_1  _077_
timestamp 1676560849
transform 1 0 4800 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _078_
timestamp 1676630787
transform 1 0 3072 0 -1 9072
box -48 -56 432 834
use sg13g2_xor2_1  _079_
timestamp 1677581577
transform 1 0 4608 0 1 9072
box -48 -56 816 834
use sg13g2_o21ai_1  _080_
timestamp 1685182643
transform 1 0 5472 0 -1 10584
box -48 -56 538 834
use sg13g2_xnor2_1  _081_
timestamp 1677520200
transform -1 0 5376 0 -1 7560
box -48 -56 816 834
use sg13g2_nand2_1  _082_
timestamp 1676560849
transform -1 0 10560 0 -1 10584
box -48 -56 432 834
use sg13g2_nand2_1  _083_
timestamp 1676560849
transform -1 0 8736 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _084_
timestamp 1676630787
transform 1 0 10944 0 -1 9072
box -48 -56 432 834
use sg13g2_xor2_1  _085_
timestamp 1677581577
transform -1 0 10560 0 -1 7560
box -48 -56 816 834
use sg13g2_o21ai_1  _086_
timestamp 1685182643
transform 1 0 8736 0 -1 9072
box -48 -56 538 834
use sg13g2_xnor2_1  _087_
timestamp 1677520200
transform 1 0 7584 0 1 7560
box -48 -56 816 834
use sg13g2_nand2_1  _088_
timestamp 1676560849
transform 1 0 9504 0 -1 12096
box -48 -56 432 834
use sg13g2_nand2_1  _089_
timestamp 1676560849
transform -1 0 7296 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _090_
timestamp 1676630787
transform 1 0 7488 0 1 10584
box -48 -56 432 834
use sg13g2_xor2_1  _091_
timestamp 1677581577
transform -1 0 8640 0 1 10584
box -48 -56 816 834
use sg13g2_o21ai_1  _092_
timestamp 1685182643
transform 1 0 8064 0 1 9072
box -48 -56 538 834
use sg13g2_xnor2_1  _093_
timestamp 1677520200
transform 1 0 7296 0 -1 10584
box -48 -56 816 834
use sg13g2_nand2_1  _094_
timestamp 1676560849
transform 1 0 4800 0 1 12096
box -48 -56 432 834
use sg13g2_nand2_1  _095_
timestamp 1676560849
transform 1 0 4224 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _096_
timestamp 1676630787
transform 1 0 3072 0 -1 12096
box -48 -56 432 834
use sg13g2_xor2_1  _097_
timestamp 1677581577
transform 1 0 3168 0 1 12096
box -48 -56 816 834
use sg13g2_o21ai_1  _098_
timestamp 1685182643
transform -1 0 5472 0 -1 10584
box -48 -56 538 834
use sg13g2_xnor2_1  _099_
timestamp 1677520200
transform 1 0 5184 0 1 10584
box -48 -56 816 834
use sg13g2_inv_1  _100_
timestamp 1676386529
transform 1 0 6048 0 1 4536
box -48 -56 336 834
use sg13g2_inv_1  _101_
timestamp 1676386529
transform -1 0 2304 0 -1 12096
box -48 -56 336 834
use sg13g2_inv_1  _102_
timestamp 1676386529
transform 1 0 1632 0 -1 9072
box -48 -56 336 834
use sg13g2_inv_1  _103_
timestamp 1676386529
transform -1 0 6336 0 -1 6048
box -48 -56 336 834
use sg13g2_inv_1  _104_
timestamp 1676386529
transform -1 0 3360 0 1 3024
box -48 -56 336 834
use sg13g2_inv_1  _105_
timestamp 1676386529
transform 1 0 4224 0 -1 9072
box -48 -56 336 834
use sg13g2_inv_1  _106_
timestamp 1676386529
transform -1 0 2208 0 -1 6048
box -48 -56 336 834
use sg13g2_inv_1  _107_
timestamp 1676386529
transform -1 0 1440 0 -1 7560
box -48 -56 336 834
use sg13g2_inv_1  _108_
timestamp 1676386529
transform -1 0 6240 0 -1 10584
box -48 -56 336 834
use sg13g2_inv_1  _109_
timestamp 1676386529
transform 1 0 5184 0 1 7560
box -48 -56 336 834
use sg13g2_inv_1  _110_
timestamp 1676386529
transform 1 0 8160 0 -1 9072
box -48 -56 336 834
use sg13g2_inv_1  _111_
timestamp 1676386529
transform 1 0 7776 0 1 9072
box -48 -56 336 834
use sg13g2_inv_1  _112_
timestamp 1676386529
transform 1 0 8448 0 -1 9072
box -48 -56 336 834
use sg13g2_inv_1  _113_
timestamp 1676386529
transform 1 0 6240 0 1 12096
box -48 -56 336 834
use sg13g2_inv_1  _114_
timestamp 1676386529
transform 1 0 2784 0 -1 12096
box -48 -56 336 834
use sg13g2_dfrbpq_1  _115_
timestamp 1746542328
transform 1 0 8736 0 -1 6048
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _116_
timestamp 1746542328
transform 1 0 7008 0 -1 4536
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _117_
timestamp 1746542328
transform 1 0 1536 0 1 10584
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _118_
timestamp 1746542328
transform 1 0 1536 0 1 9072
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _119_
timestamp 1746542328
transform 1 0 5376 0 1 3024
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _120_
timestamp 1746542328
transform 1 0 2592 0 -1 4536
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _121_
timestamp 1746542328
transform 1 0 4608 0 1 6048
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _122_
timestamp 1746542328
transform 1 0 1152 0 1 6048
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _123_
timestamp 1746542328
transform -1 0 3936 0 1 7560
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _124_
timestamp 1746542328
transform 1 0 5376 0 -1 9072
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _125_
timestamp 1746542328
transform -1 0 9312 0 -1 7560
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _126_
timestamp 1746542328
transform 1 0 8832 0 1 7560
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _127_
timestamp 1746542328
transform 1 0 8544 0 1 9072
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _128_
timestamp 1746542328
transform 1 0 8640 0 1 10584
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _129_
timestamp 1746542328
transform 1 0 6048 0 -1 12096
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _130_
timestamp 1746542328
transform 1 0 3456 0 -1 12096
box -48 -56 2640 834
use sg13g2_buf_8  clkbuf_0_clk
timestamp 1676454965
transform -1 0 7584 0 1 7560
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_2_0__f_clk
timestamp 1676454965
transform -1 0 5184 0 -1 6048
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_2_1__f_clk
timestamp 1676454965
transform 1 0 9312 0 1 6048
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_2_2__f_clk
timestamp 1676454965
transform -1 0 4128 0 -1 10584
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_2_3__f_clk
timestamp 1676454965
transform 1 0 8928 0 -1 10584
box -48 -56 1296 834
use sg13g2_buf_8  fanout1
timestamp 1676454965
transform 1 0 5376 0 -1 7560
box -48 -56 1296 834
use sg13g2_buf_8  fanout2
timestamp 1676454965
transform 1 0 6240 0 1 10584
box -48 -56 1296 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679585382
transform 1 0 1152 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679585382
transform 1 0 1824 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_14
timestamp 1679581501
transform 1 0 2496 0 1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_18
timestamp 1677583704
transform 1 0 2880 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_23
timestamp 1679585382
transform 1 0 3360 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_30
timestamp 1679585382
transform 1 0 4032 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_37
timestamp 1677583704
transform 1 0 4704 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_39
timestamp 1677583258
transform 1 0 4896 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679585382
transform 1 0 9216 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679585382
transform 1 0 9888 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679585382
transform 1 0 10560 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_105
timestamp 1677583704
transform 1 0 11232 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679585382
transform 1 0 1152 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679585382
transform 1 0 1824 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_14
timestamp 1677583258
transform 1 0 2496 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_50
timestamp 1677583704
transform 1 0 5952 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_88
timestamp 1679585382
transform 1 0 9600 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_95
timestamp 1679585382
transform 1 0 10272 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_102
timestamp 1679581501
transform 1 0 10944 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_106
timestamp 1677583258
transform 1 0 11328 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679585382
transform 1 0 1152 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679585382
transform 1 0 1824 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_14
timestamp 1677583704
transform 1 0 2496 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_71
timestamp 1677583704
transform 1 0 7968 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_73
timestamp 1677583258
transform 1 0 8160 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_83
timestamp 1679585382
transform 1 0 9120 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_90
timestamp 1679585382
transform 1 0 9792 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_97
timestamp 1679581501
transform 1 0 10464 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_101
timestamp 1677583704
transform 1 0 10848 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_11
timestamp 1677583704
transform 1 0 2208 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_106
timestamp 1677583258
transform 1 0 11328 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_63
timestamp 1677583258
transform 1 0 7200 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_76
timestamp 1679585382
transform 1 0 8448 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_83
timestamp 1677583704
transform 1 0 9120 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_98
timestamp 1677583258
transform 1 0 10560 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_25
timestamp 1677583704
transform 1 0 3552 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_57
timestamp 1677583258
transform 1 0 6624 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_85
timestamp 1679581501
transform 1 0 9312 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_89
timestamp 1677583258
transform 1 0 9696 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_0
timestamp 1677583704
transform 1 0 1152 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_79
timestamp 1677583258
transform 1 0 8736 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_0
timestamp 1679581501
transform 1 0 1152 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_4
timestamp 1677583258
transform 1 0 1536 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_13
timestamp 1677583704
transform 1 0 2400 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_15
timestamp 1677583258
transform 1 0 2592 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_71
timestamp 1677583704
transform 1 0 7968 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_106
timestamp 1677583258
transform 1 0 11328 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_31
timestamp 1677583258
transform 1 0 4128 0 1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_44
timestamp 1677583258
transform 1 0 5376 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_67
timestamp 1677583704
transform 1 0 7584 0 1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_104
timestamp 1677583704
transform 1 0 11136 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_106
timestamp 1677583258
transform 1 0 11328 0 1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_0
timestamp 1677583258
transform 1 0 1152 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_53
timestamp 1679585382
transform 1 0 6240 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_0
timestamp 1679581501
transform 1 0 1152 0 1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_31
timestamp 1677583704
transform 1 0 4128 0 1 10584
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_50
timestamp 1677583704
transform 1 0 5952 0 1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_52
timestamp 1677583258
transform 1 0 6144 0 1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_105
timestamp 1677583704
transform 1 0 11232 0 1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_12
timestamp 1679581501
transform 1 0 2304 0 -1 12096
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_16
timestamp 1677583258
transform 1 0 2688 0 -1 12096
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_100
timestamp 1679585382
transform 1 0 10752 0 -1 12096
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_0
timestamp 1679585382
transform 1 0 1152 0 1 12096
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_7
timestamp 1679585382
transform 1 0 1824 0 1 12096
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_14
timestamp 1677583704
transform 1 0 2496 0 1 12096
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_16
timestamp 1677583258
transform 1 0 2688 0 1 12096
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_42
timestamp 1677583258
transform 1 0 5184 0 1 12096
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_52
timestamp 1677583258
transform 1 0 6144 0 1 12096
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_56
timestamp 1679585382
transform 1 0 6528 0 1 12096
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_67
timestamp 1679585382
transform 1 0 7584 0 1 12096
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_74
timestamp 1679581501
transform 1 0 8256 0 1 12096
box -48 -56 432 834
use sg13g2_decap_8  FILLER_12_87
timestamp 1679585382
transform 1 0 9504 0 1 12096
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_94
timestamp 1679585382
transform 1 0 10176 0 1 12096
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_101
timestamp 1679581501
transform 1 0 10848 0 1 12096
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_105
timestamp 1677583704
transform 1 0 11232 0 1 12096
box -48 -56 240 834
use sg13g2_dlygate4sd3_1  hold1
timestamp 1677675658
transform -1 0 2880 0 -1 10584
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold2
timestamp 1677675658
transform -1 0 9120 0 1 4536
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold3
timestamp 1677675658
transform -1 0 7968 0 1 4536
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold4
timestamp 1677675658
transform -1 0 8064 0 -1 6048
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold5
timestamp 1677675658
transform -1 0 11424 0 -1 10584
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold6
timestamp 1677675658
transform -1 0 10944 0 -1 9072
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold7
timestamp 1677675658
transform -1 0 10080 0 -1 9072
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold8
timestamp 1677675658
transform -1 0 7584 0 1 9072
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold9
timestamp 1677675658
transform -1 0 6336 0 1 7560
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold10
timestamp 1677675658
transform -1 0 6336 0 1 9072
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold11
timestamp 1677675658
transform 1 0 3744 0 1 6048
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold12
timestamp 1677675658
transform -1 0 4608 0 -1 7560
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold13
timestamp 1677675658
transform -1 0 3072 0 -1 7560
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold14
timestamp 1677675658
transform 1 0 4128 0 -1 10584
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold15
timestamp 1677675658
transform 1 0 4320 0 1 10584
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold16
timestamp 1677675658
transform -1 0 4800 0 1 12096
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold17
timestamp 1677675658
transform 1 0 8640 0 1 12096
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold18
timestamp 1677675658
transform -1 0 9504 0 -1 12096
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold19
timestamp 1677675658
transform 1 0 8064 0 -1 10584
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold20
timestamp 1677675658
transform 1 0 5184 0 1 4536
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold21
timestamp 1677675658
transform -1 0 6048 0 -1 6048
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold22
timestamp 1677675658
transform -1 0 4416 0 1 4536
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold23
timestamp 1677675658
transform -1 0 4800 0 1 7560
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold24
timestamp 1677675658
transform -1 0 10752 0 -1 12096
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold25
timestamp 1677675658
transform -1 0 8832 0 1 3024
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold26
timestamp 1677675658
transform -1 0 6144 0 1 12096
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold27
timestamp 1677675658
transform -1 0 7200 0 -1 6048
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold28
timestamp 1677675658
transform -1 0 11424 0 -1 7560
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold29
timestamp 1677675658
transform 1 0 4512 0 -1 9072
box -48 -56 912 834
use sg13g2_buf_1  input1
timestamp 1676385511
transform 1 0 1632 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676385511
transform -1 0 11424 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676385511
transform -1 0 9216 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676385511
transform 1 0 1536 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676385511
transform 1 0 1152 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input6
timestamp 1676385511
transform -1 0 11424 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  input7
timestamp 1676385511
transform -1 0 7584 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  input8
timestamp 1676385511
transform 1 0 2784 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  input9
timestamp 1676385511
transform 1 0 1152 0 1 9072
box -48 -56 432 834
use sg13g2_buf_2  input10
timestamp 1676385467
transform -1 0 1632 0 -1 12096
box -48 -56 528 834
use sg13g2_buf_1  output11
timestamp 1676385511
transform 1 0 10656 0 1 6048
box -48 -56 432 834
<< labels >>
flabel metal6 s 4892 2898 5332 12896 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 1108 6764 11468 7204 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3652 2980 4092 12978 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 1108 5524 11468 5964 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 12504 4244 12584 4324 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 12504 7436 12584 7516 0 FreeSans 320 0 0 0 p
port 3 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 rst
port 4 nsew signal input
flabel metal3 s 12504 6260 12584 6340 0 FreeSans 320 0 0 0 x[0]
port 5 nsew signal input
flabel metal2 s 6968 0 7048 80 0 FreeSans 320 0 0 0 x[1]
port 6 nsew signal input
flabel metal3 s 0 5756 80 5836 0 FreeSans 320 0 0 0 x[2]
port 7 nsew signal input
flabel metal3 s 0 6932 80 7012 0 FreeSans 320 0 0 0 x[3]
port 8 nsew signal input
flabel metal3 s 12504 8780 12584 8860 0 FreeSans 320 0 0 0 x[4]
port 9 nsew signal input
flabel metal2 s 7160 16248 7240 16328 0 FreeSans 320 0 0 0 x[5]
port 10 nsew signal input
flabel metal2 s 4088 16248 4168 16328 0 FreeSans 320 0 0 0 x[6]
port 11 nsew signal input
flabel metal3 s 0 9116 80 9196 0 FreeSans 320 0 0 0 x[7]
port 12 nsew signal input
flabel metal3 s 0 11300 80 11380 0 FreeSans 320 0 0 0 y
port 13 nsew signal input
rlabel metal1 6288 12096 6288 12096 0 VGND
rlabel metal1 6288 12852 6288 12852 0 VPWR
rlabel metal2 6624 5040 6624 5040 0 _000_
rlabel metal3 3888 4872 3888 4872 0 _001_
rlabel metal2 2976 7308 2976 7308 0 _002_
rlabel metal2 6240 9912 6240 9912 0 _003_
rlabel metal3 9552 8736 9552 8736 0 _004_
rlabel metal2 8448 9828 8448 9828 0 _005_
rlabel metal2 4704 11886 4704 11886 0 _006_
rlabel metal2 1344 10626 1344 10626 0 _007_
rlabel metal2 1920 8904 1920 8904 0 _008_
rlabel metal3 8736 5712 8736 5712 0 _009_
rlabel metal2 7488 4452 7488 4452 0 _010_
rlabel metal2 2112 11424 2112 11424 0 _011_
rlabel metal2 1968 8736 1968 8736 0 _012_
rlabel metal2 5952 3360 5952 3360 0 _013_
rlabel metal2 3120 3612 3120 3612 0 _014_
rlabel metal2 5088 6888 5088 6888 0 _015_
rlabel metal2 1872 5712 1872 5712 0 _016_
rlabel metal2 1248 7476 1248 7476 0 _017_
rlabel metal2 5856 9366 5856 9366 0 _018_
rlabel metal2 8832 7392 8832 7392 0 _019_
rlabel metal3 8832 7896 8832 7896 0 _020_
rlabel metal2 9024 9324 9024 9324 0 _021_
rlabel metal2 8688 8820 8688 8820 0 _022_
rlabel metal2 6480 11760 6480 11760 0 _023_
rlabel metal2 3936 11718 3936 11718 0 _024_
rlabel metal3 4320 10164 4320 10164 0 _025_
rlabel metal3 4656 12264 4656 12264 0 _026_
rlabel metal2 6336 4326 6336 4326 0 _027_
rlabel metal2 7488 5922 7488 5922 0 _028_
rlabel metal2 6816 4830 6816 4830 0 _029_
rlabel metal2 6912 5334 6912 5334 0 _030_
rlabel metal2 2208 8778 2208 8778 0 _031_
rlabel metal2 5952 5670 5952 5670 0 _032_
rlabel metal3 4704 4872 4704 4872 0 _033_
rlabel metal2 3264 4788 3264 4788 0 _034_
rlabel metal2 5328 4284 5328 4284 0 _035_
rlabel metal3 4512 7266 4512 7266 0 _036_
rlabel metal3 3072 5712 3072 5712 0 _037_
rlabel metal3 3264 7098 3264 7098 0 _038_
rlabel metal2 3456 6258 3456 6258 0 _039_
rlabel metal2 6240 8232 6240 8232 0 _040_
rlabel metal2 5616 9408 5616 9408 0 _041_
rlabel metal3 4608 8820 4608 8820 0 _042_
rlabel metal2 4848 7224 4848 7224 0 _043_
rlabel metal2 10704 8736 10704 8736 0 _044_
rlabel metal2 8640 8148 8640 8148 0 _045_
rlabel metal2 8928 8778 8928 8778 0 _046_
rlabel metal2 9984 7518 9984 7518 0 _047_
rlabel metal2 9408 11676 9408 11676 0 _048_
rlabel metal2 7680 10080 7680 10080 0 _049_
rlabel metal2 8256 9744 8256 9744 0 _050_
rlabel metal2 7776 10500 7776 10500 0 _051_
rlabel metal3 4704 12348 4704 12348 0 _052_
rlabel metal3 4896 10248 4896 10248 0 _053_
rlabel metal2 7296 7014 7296 7014 0 clk
rlabel metal3 5328 7896 5328 7896 0 clknet_0_clk
rlabel metal2 3936 4116 3936 4116 0 clknet_2_0__leaf_clk
rlabel metal2 10080 6006 10080 6006 0 clknet_2_1__leaf_clk
rlabel metal3 4128 11760 4128 11760 0 clknet_2_2__leaf_clk
rlabel metal3 7056 10080 7056 10080 0 clknet_2_3__leaf_clk
rlabel metal2 8832 6132 8832 6132 0 csa0.hsum2
rlabel metal2 9504 4620 9504 4620 0 csa0.sc
rlabel metal2 8736 3864 8736 3864 0 csa0.y
rlabel metal2 5520 3360 5520 3360 0 genblk1\[1\].csa.hsum2
rlabel metal3 5232 4368 5232 4368 0 genblk1\[1\].csa.sc
rlabel metal2 7104 5964 7104 5964 0 genblk1\[1\].csa.y
rlabel metal3 4272 5880 4272 5880 0 genblk1\[2\].csa.hsum2
rlabel metal2 3840 6426 3840 6426 0 genblk1\[2\].csa.sc
rlabel metal2 1920 7476 1920 7476 0 genblk1\[2\].csa.y
rlabel metal3 4272 7392 4272 7392 0 genblk1\[3\].csa.hsum2
rlabel metal2 7872 8736 7872 8736 0 genblk1\[3\].csa.sc
rlabel metal2 6624 8400 6624 8400 0 genblk1\[3\].csa.y
rlabel metal2 9216 7518 9216 7518 0 genblk1\[4\].csa.hsum2
rlabel metal2 11328 9198 11328 9198 0 genblk1\[4\].csa.sc
rlabel metal2 11232 7980 11232 7980 0 genblk1\[4\].csa.y
rlabel metal3 8304 9408 8304 9408 0 genblk1\[5\].csa.hsum2
rlabel metal2 9792 11718 9792 11718 0 genblk1\[5\].csa.sc
rlabel metal2 8544 12180 8544 12180 0 genblk1\[5\].csa.y
rlabel metal2 6144 11550 6144 11550 0 genblk1\[6\].csa.hsum2
rlabel metal2 5088 12516 5088 12516 0 genblk1\[6\].csa.sc
rlabel metal2 4224 10500 4224 10500 0 genblk1\[6\].csa.y
rlabel metal2 6144 4284 6144 4284 0 net1
rlabel metal3 3696 11928 3696 11928 0 net10
rlabel metal2 1440 8988 1440 8988 0 net11
rlabel metal2 1440 11550 1440 11550 0 net12
rlabel metal2 11232 6174 11232 6174 0 net13
rlabel metal2 2208 10080 2208 10080 0 net14
rlabel metal3 8496 5040 8496 5040 0 net15
rlabel metal2 6720 4326 6720 4326 0 net16
rlabel metal2 7200 4200 7200 4200 0 net17
rlabel metal2 11040 8652 11040 8652 0 net18
rlabel metal2 9024 8694 9024 8694 0 net19
rlabel metal2 2304 11760 2304 11760 0 net2
rlabel metal2 8928 8190 8928 8190 0 net20
rlabel metal3 3936 9408 3936 9408 0 net21
rlabel metal2 5664 8148 5664 8148 0 net22
rlabel metal2 5520 8820 5520 8820 0 net23
rlabel metal2 2112 7140 2112 7140 0 net24
rlabel metal3 3600 7224 3600 7224 0 net25
rlabel metal3 1776 6384 1776 6384 0 net26
rlabel metal2 4896 12474 4896 12474 0 net27
rlabel metal2 5184 10332 5184 10332 0 net28
rlabel metal3 3792 11844 3792 11844 0 net29
rlabel metal4 1920 12180 1920 12180 0 net3
rlabel metal3 8928 11760 8928 11760 0 net30
rlabel metal2 8736 11424 8736 11424 0 net31
rlabel metal2 8784 10416 8784 10416 0 net32
rlabel metal2 3024 4872 3024 4872 0 net33
rlabel metal2 3360 4956 3360 4956 0 net34
rlabel metal2 2688 4368 2688 4368 0 net35
rlabel metal2 4080 8148 4080 8148 0 net36
rlabel metal3 9264 11508 9264 11508 0 net37
rlabel metal2 8064 4242 8064 4242 0 net38
rlabel metal3 4320 12432 4320 12432 0 net39
rlabel metal2 11136 5670 11136 5670 0 net4
rlabel metal2 5472 4830 5472 4830 0 net40
rlabel metal3 10368 7224 10368 7224 0 net41
rlabel metal2 5328 8904 5328 8904 0 net42
rlabel metal3 7104 3360 7104 3360 0 net5
rlabel metal2 2496 5796 2496 5796 0 net6
rlabel metal2 1440 5922 1440 5922 0 net7
rlabel metal2 11136 7308 11136 7308 0 net8
rlabel metal2 7296 11802 7296 11802 0 net9
rlabel metal2 10944 7056 10944 7056 0 p
rlabel metal3 894 11508 894 11508 0 rst
rlabel metal3 4080 9660 4080 9660 0 tcmp.z
rlabel metal3 11926 6300 11926 6300 0 x[0]
rlabel metal2 7008 660 7008 660 0 x[1]
rlabel metal3 846 5796 846 5796 0 x[2]
rlabel metal3 606 6972 606 6972 0 x[3]
rlabel metal3 11974 8820 11974 8820 0 x[4]
rlabel metal2 7200 14396 7200 14396 0 x[5]
rlabel metal2 4128 15068 4128 15068 0 x[6]
rlabel metal3 654 9156 654 9156 0 x[7]
rlabel metal2 1248 11550 1248 11550 0 y
<< properties >>
string FIXED_BBOX 0 0 12584 16328
<< end >>
