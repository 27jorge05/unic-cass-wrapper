* Extracted by KLayout with SG13G2 LVS runset on : 15/01/2026 11:02

.SUBCKT user_project_wrapper VDD VSS ui_PAD[9] ui_PAD[10] ui_PAD[11] ui_PAD[12]
+ ui_PAD[13] ui_PAD[14] ui_PAD[15] analog_io_0 io_clock_PAD IOVDD IOVSS
+ ui_PAD[0] uo_PAD[0] ui_PAD[1] uo_PAD[1] ui_PAD[2] uo_PAD[2] ui_PAD[3]
+ uo_PAD[3] ui_PAD[4] uo_PAD[4] ui_PAD[5] uo_PAD[5] ui_PAD[6] uo_PAD[6]
+ ui_PAD[7] uo_PAD[7] ui_PAD[8] uo_PAD[8] uo_PAD[9] uo_PAD[10] uo_PAD[11]
+ uo_PAD[12] uo_PAD[13] uo_PAD[14] uo_PAD[15] analog_io_1 io_reset_PAD
X$1 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$2 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Corner
X$3 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler1000
X$4 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$5 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler200
X$6 \$1 VDD IOVSS IOVSS VSS sg13g2_IOPadVdd
X$8 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$9 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$10 \$1 VSS IOVSS IOVSS IOVDD sg13g2_IOPadVss
X$12 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$13 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$14 \$1 ui_PAD[9] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$16 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$17 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$18 \$1 ui_PAD[10] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$20 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$21 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$22 \$1 ui_PAD[11] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$24 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$25 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$26 \$1 ui_PAD[12] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$28 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$29 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$30 \$1 ui_PAD[13] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$32 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$33 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$34 \$1 ui_PAD[14] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$36 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$37 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$38 \$1 ui_PAD[15] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$40 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$41 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$42 \$1 analog_io_0 IOVSS IOVDD IOVDD VSS sg13g2_IOPadAnalog
X$44 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$45 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$46 \$1 io_clock_PAD IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$48 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$49 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$50 \$1 IOVDD IOVSS IOVSS VSS sg13g2_IOPadIOVdd
X$52 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$53 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$54 \$1 IOVSS IOVDD VSS sg13g2_IOPadIOVss
X$56 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$57 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler1000
X$58 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$59 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler200
X$60 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Corner
X$61 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$62 \$1 VDD IOVSS IOVSS VSS sg13g2_IOPadVdd
X$64 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$65 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$66 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler200
X$67 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$68 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler1000
X$69 \$1 VSS IOVSS IOVSS IOVDD sg13g2_IOPadVss
X$71 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$72 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$73 \$1 ui_PAD[0] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$75 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$76 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$77 \$1 ui_PAD[1] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$79 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$80 \$1 ui_PAD[4] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$82 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$83 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$84 \$1 ui_PAD[3] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$86 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$87 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$88 \$1 ui_PAD[2] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$90 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$91 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$92 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler1000
X$93 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$94 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler200
X$95 \$1 VDD IOVSS IOVSS VSS sg13g2_IOPadVdd
X$96 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$97 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$98 \$1 uo_PAD[2] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$99 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$100 \$1 uo_PAD[3] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$101 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$102 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$103 \$1 uo_PAD[4] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$104 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$105 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$106 \$1 uo_PAD[1] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$107 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$108 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$109 \$1 uo_PAD[0] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$110 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$111 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$112 \$1 VSS IOVSS IOVSS IOVDD sg13g2_IOPadVss
X$113 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$121 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$122 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$123 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$124 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$125 \$1 ui_PAD[5] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$127 \$1 uo_PAD[5] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$129 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$130 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$131 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$132 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$133 \$1 ui_PAD[6] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$135 \$1 uo_PAD[6] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$137 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$138 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$139 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$140 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$141 \$1 ui_PAD[7] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$143 \$1 uo_PAD[7] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$145 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$146 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$147 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$148 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$149 \$1 ui_PAD[8] IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$151 \$1 uo_PAD[8] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$153 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$154 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$155 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$156 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$157 \$1 IOVDD IOVSS IOVSS VSS sg13g2_IOPadIOVdd
X$159 \$1 IOVDD IOVSS IOVSS VSS sg13g2_IOPadIOVdd
X$161 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$162 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$163 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$164 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$165 \$1 IOVSS IOVDD VSS sg13g2_IOPadIOVss
X$167 \$1 IOVSS IOVDD VSS sg13g2_IOPadIOVss
X$169 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$170 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler1000
X$171 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$172 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler1000
X$173 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$174 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler200
X$175 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$176 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler200
X$177 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Corner
X$178 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$179 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler1000
X$180 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$181 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler200
X$182 \$1 IOVDD IOVSS IOVSS VSS sg13g2_IOPadIOVdd
X$183 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$184 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$185 \$1 IOVSS IOVDD VSS sg13g2_IOPadIOVss
X$186 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$187 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$188 \$1 uo_PAD[9] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$189 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$190 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$191 \$1 uo_PAD[10] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$192 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$193 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$194 \$1 uo_PAD[11] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$195 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$196 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$197 \$1 uo_PAD[12] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$198 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$199 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$200 \$1 uo_PAD[13] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$201 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$202 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$203 \$1 uo_PAD[14] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$204 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$205 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$206 \$1 uo_PAD[15] IOVSS IOVDD IOVDD VDD VSS sg13g2_IOPadOut30mA
X$207 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$208 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$209 \$1 analog_io_1 IOVSS IOVDD IOVDD VSS sg13g2_IOPadAnalog
X$210 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$211 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$212 \$1 io_reset_PAD IOVSS IOVSS IOVDD VDD VSS sg13g2_IOPadIn
X$213 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$214 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$215 \$1 IOVDD IOVSS IOVSS VSS sg13g2_IOPadIOVdd
X$216 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$217 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$218 \$1 IOVSS IOVDD VSS sg13g2_IOPadIOVss
X$219 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler4000
X$220 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler1000
X$221 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler400
X$222 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Filler200
X$223 \$1 IOVSS IOVSS IOVSS VSS sg13g2_Corner
.ENDS user_project_wrapper

.SUBCKT sg13g2_IOPadVss \$1 vss iovss iovss$1 iovdd
R$1 \$1 iovss$1 ptap1 A=5407.1p P=703.48u
R$2 \$1 vss ptap1 A=24p P=160.6u
D$3 vss iovdd dpantenna A=35.0028p P=58.08u m=2
D$5 \$1 vss dantenna A=35.0028p P=58.08u m=2
R$7 \$1 iovss ptap1 A=141.2964p P=221.76u
.ENDS sg13g2_IOPadVss

.SUBCKT sg13g2_IOPadVdd \$1 vdd iovss iovss$1 vss
R$1 \$1 iovss$1 ptap1 A=2051.93485p P=727.53u
R$2 \$1 vss ptap1 A=24p P=160.6u
M$3 iovss$1 vdd iovss$1 \$1 sg13_hv_nmos L=9.5u W=126u AS=26.64p AD=23.94p
+ PS=149.92u PD=131.32u
M$10 iovss$1 vdd \$10 \$1 sg13_hv_nmos L=0.5u W=108u AS=20.52p AD=23.22p
+ PS=112.56u PD=131.16u
M$29 vdd vdd \$10 vdd sg13_hv_pmos L=0.5u W=350u AS=67.55p AD=67.55p PS=376.3u
+ PD=376.3u
M$79 iovss \$10 vdd \$1 sg13_hv_nmos L=0.6u W=756.8u AS=344.608p AD=349.36p
+ PS=931.04u PD=933.2u
D$251 \$1 \$10 dantenna A=0.2304p P=1.92u m=1
R$252 \$1 iovss ptap1 A=65.6472p P=386.16u
.ENDS sg13g2_IOPadVdd

.SUBCKT sg13g2_IOPadAnalog \$1 pad|padres iovss iovdd iovdd$1 vss
R$1 \$1 iovss ptap1 A=4580.0452p P=1715.26u
R$2 \$1 vss ptap1 A=23.85p P=159.6u
M$6 iovdd \$I15 pad|padres iovdd sg13_hv_pmos L=0.6u W=266.4u AS=123.21p
+ AD=123.21p PS=316.72u PD=316.72u
R$46 iovdd \$I15 rppd w=0.5u l=12.9u ps=0 b=0 m=1
M$47 iovss \$I16 pad|padres \$1 sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p
+ PS=110.9u PD=110.9u
R$67 iovss \$I16 rppd w=0.5u l=3.54u ps=0 b=0 m=1
D$69 pad|padres iovdd dpantenna A=35.0028p P=58.08u m=2
D$71 \$1 pad|padres dantenna A=35.0028p P=58.08u m=2
D$74 \$1 pad|padres dantenna A=1.984p P=7.48u m=1
D$75 pad|padres iovdd$1 dpantenna A=3.1872p P=11.24u m=1
.ENDS sg13g2_IOPadAnalog

.SUBCKT sg13g2_IOPadIOVss \$1 iovss iovdd vss
R$1 \$1 iovss ptap1 A=5548.3964p P=925.24u
R$2 \$1 vss ptap1 A=24p P=160.6u
D$3 iovss iovdd dpantenna A=35.0028p P=58.08u m=2
D$5 \$1 iovss dantenna A=35.0028p P=58.08u m=2
.ENDS sg13g2_IOPadIOVss

.SUBCKT sg13g2_IOPadIOVdd \$1 iovdd iovss iovss$1 vss
R$1 \$1 iovss$1 ptap1 A=2052.0763p P=727.52u
R$2 \$1 vss ptap1 A=24p P=160.6u
M$3 iovss$1 iovdd iovss$1 \$1 sg13_hv_nmos L=9.5u W=126u AS=26.64p AD=23.94p
+ PS=149.92u PD=131.32u
M$10 iovss$1 iovdd \$7 \$1 sg13_hv_nmos L=0.5u W=108u AS=20.52p AD=23.22p
+ PS=112.56u PD=131.16u
M$29 iovdd iovdd \$7 iovdd sg13_hv_pmos L=0.5u W=350u AS=67.55p AD=67.55p
+ PS=376.3u PD=376.3u
M$79 iovss \$7 iovdd \$1 sg13_hv_nmos L=0.6u W=756.8u AS=344.608p AD=349.36p
+ PS=931.04u PD=933.2u
D$251 \$1 \$7 dantenna A=0.2304p P=1.92u m=1
R$252 \$1 iovss ptap1 A=65.6472p P=386.16u
.ENDS sg13g2_IOPadIOVdd

.SUBCKT sg13g2_Filler200 \$1 iovss iovss$1 iovss$2 vss
R$1 \$1 iovss ptap1 A=13.7536p P=50.24u
R$2 \$1 iovss$1 ptap1 A=13.4736p P=49.24u
R$3 \$1 iovss$2 ptap1 A=13.748p P=50.22u
R$4 \$1 vss ptap1 A=0.678p P=5.12u
.ENDS sg13g2_Filler200

.SUBCKT sg13g2_Filler400 \$1 iovss iovss$1 iovss$2 vss
R$1 \$1 iovss ptap1 A=38.3136p P=52.24u
R$2 \$1 iovss$1 ptap1 A=37.5336p P=51.24u
R$3 \$1 iovss$2 ptap1 A=38.298p P=52.22u
R$4 \$1 vss ptap1 A=0.672p P=5.08u
.ENDS sg13g2_Filler400

.SUBCKT sg13g2_Filler1000 \$1 iovss iovss$1 iovss$2 vss
R$1 \$1 iovss ptap1 A=110.52p P=58.12u
R$2 \$1 iovss$1 ptap1 A=108.27p P=57.12u
R$3 \$1 iovss$2 ptap1 A=110.475p P=58.1u
R$4 \$1 vss ptap1 A=1.368p P=9.72u
.ENDS sg13g2_Filler1000

.SUBCKT sg13g2_Filler4000 \$1 iovss iovss$1 iovss$2 vss
R$1 \$1 iovss ptap1 A=478.92p P=88.12u
R$2 \$1 iovss$1 ptap1 A=469.17p P=87.12u
R$3 \$1 iovss$2 ptap1 A=478.725p P=88.1u
R$4 \$1 vss ptap1 A=5.85p P=39.6u
.ENDS sg13g2_Filler4000

.SUBCKT sg13g2_Corner \$1 iovss iovss$1 iovss$2 vss
R$1 \$1 iovss ptap1 A=4546.51p P=420.331u
R$2 \$1 iovss$1 ptap1 A=3344.1864p P=326.866u
R$3 \$1 iovss$2 ptap1 A=2278.0436p P=235.225u
R$4 \$1 vss ptap1 A=13.1934p P=84.704u
.ENDS sg13g2_Corner

.SUBCKT sg13g2_IOPadOut30mA \$1 pad iovss iovdd iovdd$1 vdd vss
X$1 iovdd$1 vdd vss \$27 \$5 c2p \$1 sg13g2_GateLevelUpInv
X$3 \$1 iovss pad pad pad pad pad pad pad pad \$5 sg13g2_Clamp_N15N15D
X$5 iovdd pad pad pad pad pad pad pad pad \$27 sg13g2_Clamp_P15N15D
R$1 \$1 vss ptap1 A=24p P=160.6u
R$2 \$1 iovss ptap1 A=4555.2412p P=1175.06u
D$3 pad iovdd dpantenna A=35.0028p P=58.08u m=2
D$5 \$1 pad dantenna A=35.0028p P=58.08u m=2
.ENDS sg13g2_IOPadOut30mA

.SUBCKT sg13g2_IOPadIn \$1 pad iovss iovss$1 iovdd vdd vss
R$1 \$1 vss ptap1 A=24p P=160.6u
R$2 \$1 iovss$1 ptap1 A=5416.1304p P=746.28u
M$3 p2c \$I13 vss \$1 sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u
+ PD=6.18u
M$4 vss pad \$I13 \$1 sg13_hv_nmos L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u
+ PD=5.98u
M$5 p2c \$I13 vdd vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$6 vdd pad \$I13 vdd sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u
+ PD=9.98u
D$7 pad iovdd dpantenna A=35.0028p P=58.08u m=2
D$9 \$1 pad dantenna A=35.0028p P=58.08u m=2
R$11 \$1 iovss ptap1 A=141.2964p P=221.76u
D$12 \$1 pad dantenna A=1.984p P=7.48u m=1
D$13 pad iovdd dpantenna A=3.1872p P=11.24u m=1
.ENDS sg13g2_IOPadIn

.SUBCKT sg13g2_GateLevelUpInv iovdd vdd vss pgate ngate core \$7
X$1 iovdd ngate \$7 core vss vdd sg13g2_LevelUpInv
X$2 iovdd pgate \$7 core vss vdd sg13g2_LevelUpInv
.ENDS sg13g2_GateLevelUpInv

.SUBCKT sg13g2_Clamp_N15N15D \$2 iovss pad pad$1 pad$2 pad$3 pad$4 pad$5 pad$6
+ pad$7 gate
M$1 iovss gate pad \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.664p AD=4.004p PS=15.32u
+ PD=10.62u
M$3 iovss gate pad$1 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$5 iovss gate pad$2 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$7 iovss gate pad$3 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$9 iovss gate pad$4 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$11 iovss gate pad$5 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$13 iovss gate pad$6 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$15 iovss gate pad$7 \$2 sg13_hv_nmos L=0.6u W=4.4u AS=1.408p AD=3.256p
+ PS=5.04u PD=10.28u
D$16 \$2 gate dantenna A=0.6084p P=3.12u m=1
R$17 \$2 iovss ptap1 A=55.7736p P=328.08u
.ENDS sg13g2_Clamp_N15N15D

.SUBCKT sg13g2_Clamp_P15N15D iovdd pad pad$1 pad$2 pad$3 pad$4 pad$5 pad$6
+ pad$7 gate
M$1 iovdd gate pad iovdd sg13_hv_pmos L=0.6u W=26.64u AS=14.1192p AD=12.1212p
+ PS=44.2u PD=30.28u
M$3 iovdd gate pad$1 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p AD=12.1212p
+ PS=30.28u PD=30.28u
M$5 iovdd gate pad$2 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p AD=12.1212p
+ PS=30.28u PD=30.28u
M$7 iovdd gate pad$3 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p AD=12.1212p
+ PS=30.28u PD=30.28u
M$9 iovdd gate pad$4 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p AD=12.1212p
+ PS=30.28u PD=30.28u
M$11 iovdd gate pad$5 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p
+ AD=12.1212p PS=30.28u PD=30.28u
M$13 iovdd gate pad$6 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p
+ AD=12.1212p PS=30.28u PD=30.28u
M$15 iovdd gate pad$7 iovdd sg13_hv_pmos L=0.6u W=13.32u AS=4.2624p AD=9.8568p
+ PS=14.6u PD=29.6u
D$31 gate iovdd dpantenna A=0.6084p P=3.12u m=1
.ENDS sg13g2_Clamp_P15N15D

.SUBCKT sg13g2_LevelUpInv iovdd o \$5 i vss vdd
M$1 \$6 i vss \$5 sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u
+ PD=6.18u
M$2 vss \$4 o \$5 sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u
+ PD=4.48u
M$3 \$3 i vss \$5 sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p PS=4.48u
+ PD=2.28u
M$4 vss \$6 \$4 \$5 sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u
+ PD=4.48u
M$5 \$6 i vdd vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p PS=10.18u
+ PD=10.18u
M$6 iovdd \$4 o iovdd sg13_hv_pmos L=0.45u W=3.9u AS=1.326p AD=1.326p PS=8.48u
+ PD=8.48u
M$7 \$3 \$4 iovdd iovdd sg13_hv_pmos L=0.45u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$8 iovdd \$3 \$4 iovdd sg13_hv_pmos L=0.45u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
.ENDS sg13g2_LevelUpInv
