* NGSPICE file created from spm.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

.subckt spm VGND VPWR clk p rst x[0] x[1] x[2] x[3] x[4] x[5] x[6] x[7] y
XFILLER_12_87 VPWR VGND sg13g2_decap_8
X_062_ _008_ _031_ net14 VPWR VGND sg13g2_nand2b_1
X_114_ VPWR _024_ net2 VGND sg13g2_inv_1
X_130_ _024_ VGND VPWR net29 genblk1\[6\].csa.sc clknet_2_2__leaf_clk sg13g2_dfrbpq_1
X_113_ VPWR _023_ net3 VGND sg13g2_inv_1
X_061_ _031_ net12 net11 VPWR VGND sg13g2_nand2_1
XFILLER_0_14 VPWR VGND sg13g2_decap_4
XFILLER_6_79 VPWR VGND sg13g2_fill_1
Xhold20 genblk1\[1\].csa.sc VPWR VGND net33 sg13g2_dlygate4sd3_1
XFILLER_12_67 VPWR VGND sg13g2_decap_8
XFILLER_12_56 VPWR VGND sg13g2_decap_8
XFILLER_10_105 VPWR VGND sg13g2_fill_2
XFILLER_0_37 VPWR VGND sg13g2_fill_2
XFILLER_2_101 VPWR VGND sg13g2_fill_2
X_060_ csa0.hsum2 _028_ _030_ VPWR VGND sg13g2_xnor2_1
Xhold10 _003_ VPWR VGND net23 sg13g2_dlygate4sd3_1
X_112_ VPWR _022_ net1 VGND sg13g2_inv_1
XFILLER_1_0 VPWR VGND sg13g2_decap_8
Xhold21 _032_ VPWR VGND net34 sg13g2_dlygate4sd3_1
Xoutput11 net13 p VPWR VGND sg13g2_buf_1
X_111_ VPWR _021_ net1 VGND sg13g2_inv_1
Xhold22 _001_ VPWR VGND net35 sg13g2_dlygate4sd3_1
Xhold11 genblk1\[2\].csa.sc VPWR VGND net24 sg13g2_dlygate4sd3_1
XFILLER_12_14 VPWR VGND sg13g2_fill_2
XFILLER_0_39 VPWR VGND sg13g2_fill_1
X_110_ VPWR _020_ net1 VGND sg13g2_inv_1
Xhold23 genblk1\[2\].csa.y VPWR VGND net36 sg13g2_dlygate4sd3_1
Xhold12 _036_ VPWR VGND net25 sg13g2_dlygate4sd3_1
XFILLER_0_18 VPWR VGND sg13g2_fill_2
Xhold24 genblk1\[5\].csa.sc VPWR VGND net37 sg13g2_dlygate4sd3_1
XFILLER_1_50 VPWR VGND sg13g2_fill_2
Xhold13 _002_ VPWR VGND net26 sg13g2_dlygate4sd3_1
XFILLER_7_71 VPWR VGND sg13g2_fill_2
XFILLER_12_16 VPWR VGND sg13g2_fill_1
XFILLER_4_83 VPWR VGND sg13g2_fill_2
X_099_ genblk1\[6\].csa.hsum2 _053_ _026_ VPWR VGND sg13g2_xnor2_1
Xhold14 genblk1\[6\].csa.y VPWR VGND net27 sg13g2_dlygate4sd3_1
Xhold25 csa0.y VPWR VGND net38 sg13g2_dlygate4sd3_1
XFILLER_1_95 VPWR VGND sg13g2_decap_8
Xhold26 genblk1\[6\].csa.sc VPWR VGND net39 sg13g2_dlygate4sd3_1
XFILLER_10_50 VPWR VGND sg13g2_fill_2
X_098_ net28 VPWR _006_ VGND _053_ _025_ sg13g2_o21ai_1
Xhold15 _052_ VPWR VGND net28 sg13g2_dlygate4sd3_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_4_63 VPWR VGND sg13g2_fill_1
X_097_ net27 net39 _026_ VPWR VGND sg13g2_xor2_1
Xhold16 _006_ VPWR VGND net29 sg13g2_dlygate4sd3_1
Xhold27 genblk1\[1\].csa.y VPWR VGND net40 sg13g2_dlygate4sd3_1
Xclkbuf_2_0__f_clk clknet_0_clk clknet_2_0__leaf_clk VPWR VGND sg13g2_buf_8
Xhold17 genblk1\[5\].csa.y VPWR VGND net30 sg13g2_dlygate4sd3_1
X_096_ genblk1\[6\].csa.sc net27 _025_ VPWR VGND sg13g2_nor2_1
XFILLER_10_52 VPWR VGND sg13g2_fill_1
XFILLER_1_7 VPWR VGND sg13g2_decap_8
Xhold28 genblk1\[4\].csa.y VPWR VGND net41 sg13g2_dlygate4sd3_1
X_079_ net42 net21 _043_ VPWR VGND sg13g2_xor2_1
XFILLER_4_76 VPWR VGND sg13g2_decap_8
XFILLER_4_98 VPWR VGND sg13g2_fill_1
X_095_ _053_ net12 net10 VPWR VGND sg13g2_nand2_1
XFILLER_1_88 VPWR VGND sg13g2_decap_8
Xhold18 _048_ VPWR VGND net31 sg13g2_dlygate4sd3_1
XFILLER_10_31 VPWR VGND sg13g2_fill_2
Xhold29 genblk1\[3\].csa.y VPWR VGND net42 sg13g2_dlygate4sd3_1
X_078_ net21 genblk1\[3\].csa.y _042_ VPWR VGND sg13g2_nor2_1
XFILLER_8_104 VPWR VGND sg13g2_fill_2
X_094_ _052_ genblk1\[6\].csa.sc net27 VPWR VGND sg13g2_nand2_1
Xhold19 _005_ VPWR VGND net32 sg13g2_dlygate4sd3_1
X_129_ _023_ VGND VPWR genblk1\[6\].csa.hsum2 genblk1\[5\].csa.y clknet_2_3__leaf_clk
+ sg13g2_dfrbpq_1
X_077_ _041_ net12 net7 VPWR VGND sg13g2_nand2_1
XFILLER_12_101 VPWR VGND sg13g2_decap_4
X_093_ genblk1\[5\].csa.hsum2 _049_ _051_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_0 VPWR VGND sg13g2_fill_2
Xinput1 rst net3 VPWR VGND sg13g2_buf_1
X_076_ _040_ net21 genblk1\[3\].csa.y VPWR VGND sg13g2_nand2_1
X_128_ _022_ VGND VPWR net32 genblk1\[5\].csa.sc clknet_2_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_8_106 VPWR VGND sg13g2_fill_1
X_059_ net16 VPWR _000_ VGND _028_ _029_ sg13g2_o21ai_1
X_092_ net31 VPWR _005_ VGND _049_ _050_ sg13g2_o21ai_1
XFILLER_1_14 VPWR VGND sg13g2_fill_1
Xinput2 x[0] net4 VPWR VGND sg13g2_buf_1
X_127_ _021_ VGND VPWR genblk1\[5\].csa.hsum2 genblk1\[4\].csa.y clknet_2_3__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_7_13 VPWR VGND sg13g2_fill_2
X_058_ net38 net15 _030_ VPWR VGND sg13g2_xor2_1
XFILLER_2_90 VPWR VGND sg13g2_decap_8
X_075_ genblk1\[2\].csa.hsum2 _037_ _039_ VPWR VGND sg13g2_xnor2_1
XFILLER_1_102 VPWR VGND sg13g2_decap_4
X_091_ net30 net37 _051_ VPWR VGND sg13g2_xor2_1
Xinput3 x[1] net5 VPWR VGND sg13g2_buf_1
X_074_ net25 VPWR _002_ VGND _037_ _038_ sg13g2_o21ai_1
X_126_ _020_ VGND VPWR net20 genblk1\[4\].csa.sc clknet_2_1__leaf_clk sg13g2_dfrbpq_1
X_057_ net15 csa0.y _029_ VPWR VGND sg13g2_nor2_1
X_109_ VPWR _019_ net1 VGND sg13g2_inv_1
X_090_ genblk1\[5\].csa.sc net30 _050_ VPWR VGND sg13g2_nor2_1
Xinput4 x[2] net6 VPWR VGND sg13g2_buf_1
Xclkbuf_2_1__f_clk clknet_0_clk clknet_2_1__leaf_clk VPWR VGND sg13g2_buf_8
X_073_ net36 net24 _039_ VPWR VGND sg13g2_xor2_1
XFILLER_7_15 VPWR VGND sg13g2_fill_1
X_056_ _028_ net12 net4 VPWR VGND sg13g2_nand2_1
X_125_ _019_ VGND VPWR genblk1\[4\].csa.hsum2 genblk1\[3\].csa.y clknet_2_1__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_12_105 VPWR VGND sg13g2_fill_2
X_108_ VPWR _018_ net2 VGND sg13g2_inv_1
Xinput5 x[3] net7 VPWR VGND sg13g2_buf_1
X_072_ net24 genblk1\[2\].csa.y _038_ VPWR VGND sg13g2_nor2_1
X_124_ _018_ VGND VPWR net23 genblk1\[3\].csa.sc clknet_2_3__leaf_clk sg13g2_dfrbpq_1
X_055_ _027_ net15 csa0.y VPWR VGND sg13g2_nand2_1
XFILLER_2_71 VPWR VGND sg13g2_fill_2
XFILLER_12_0 VPWR VGND sg13g2_decap_8
X_107_ VPWR _017_ net2 VGND sg13g2_inv_1
XFILLER_2_83 VPWR VGND sg13g2_decap_8
X_071_ _037_ net12 net6 VPWR VGND sg13g2_nand2_1
Xinput6 x[4] net8 VPWR VGND sg13g2_buf_1
X_106_ VPWR _016_ net2 VGND sg13g2_inv_1
X_054_ VPWR _009_ net1 VGND sg13g2_inv_1
X_123_ _017_ VGND VPWR genblk1\[3\].csa.hsum2 genblk1\[2\].csa.y clknet_2_2__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_1_106 VPWR VGND sg13g2_fill_1
Xinput7 x[5] net9 VPWR VGND sg13g2_buf_1
X_070_ _036_ net24 genblk1\[2\].csa.y VPWR VGND sg13g2_nand2_1
Xinput10 y net12 VPWR VGND sg13g2_buf_2
XFILLER_2_0 VPWR VGND sg13g2_decap_8
XFILLER_2_73 VPWR VGND sg13g2_fill_1
X_122_ _016_ VGND VPWR net26 genblk1\[2\].csa.sc clknet_2_0__leaf_clk sg13g2_dfrbpq_1
X_105_ VPWR _015_ net2 VGND sg13g2_inv_1
Xinput8 x[6] net10 VPWR VGND sg13g2_buf_1
X_104_ VPWR _014_ net1 VGND sg13g2_inv_1
X_121_ _015_ VGND VPWR genblk1\[2\].csa.hsum2 genblk1\[1\].csa.y clknet_2_0__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_10_0 VPWR VGND sg13g2_decap_4
Xinput9 x[7] net11 VPWR VGND sg13g2_buf_1
XFILLER_5_85 VPWR VGND sg13g2_decap_4
X_120_ _014_ VGND VPWR net35 genblk1\[1\].csa.sc clknet_2_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_2_97 VPWR VGND sg13g2_decap_4
X_103_ VPWR _013_ net1 VGND sg13g2_inv_1
Xhold1 tcmp.z VPWR VGND net14 sg13g2_dlygate4sd3_1
XFILLER_11_100 VPWR VGND sg13g2_decap_8
Xclkbuf_2_2__f_clk clknet_0_clk clknet_2_2__leaf_clk VPWR VGND sg13g2_buf_8
X_102_ VPWR _012_ net2 VGND sg13g2_inv_1
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_8_31 VPWR VGND sg13g2_fill_1
Xhold2 csa0.sc VPWR VGND net15 sg13g2_dlygate4sd3_1
X_101_ VPWR _011_ net2 VGND sg13g2_inv_1
Xhold3 _027_ VPWR VGND net16 sg13g2_dlygate4sd3_1
XFILLER_7_106 VPWR VGND sg13g2_fill_1
X_100_ VPWR _010_ net1 VGND sg13g2_inv_1
XFILLER_12_7 VPWR VGND sg13g2_decap_8
XFILLER_8_44 VPWR VGND sg13g2_fill_1
Xhold4 _000_ VPWR VGND net17 sg13g2_dlygate4sd3_1
XFILLER_5_89 VPWR VGND sg13g2_fill_1
XFILLER_8_67 VPWR VGND sg13g2_fill_2
Xhold5 genblk1\[4\].csa.sc VPWR VGND net18 sg13g2_dlygate4sd3_1
XFILLER_5_57 VPWR VGND sg13g2_fill_1
XFILLER_11_12 VPWR VGND sg13g2_decap_4
XFILLER_9_0 VPWR VGND sg13g2_fill_1
XFILLER_2_14 VPWR VGND sg13g2_fill_2
XFILLER_2_7 VPWR VGND sg13g2_decap_8
X_089_ _049_ net12 net9 VPWR VGND sg13g2_nand2_1
Xhold6 _044_ VPWR VGND net19 sg13g2_dlygate4sd3_1
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_5_25 VPWR VGND sg13g2_fill_2
X_088_ _048_ genblk1\[5\].csa.sc net30 VPWR VGND sg13g2_nand2_1
Xhold7 _004_ VPWR VGND net20 sg13g2_dlygate4sd3_1
Xhold8 genblk1\[3\].csa.sc VPWR VGND net21 sg13g2_dlygate4sd3_1
X_087_ genblk1\[4\].csa.hsum2 _045_ _047_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_2_3__f_clk clknet_0_clk clknet_2_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_0_105 VPWR VGND sg13g2_fill_2
X_086_ net19 VPWR _004_ VGND _045_ _046_ sg13g2_o21ai_1
XFILLER_7_0 VPWR VGND sg13g2_decap_4
XFILLER_0_7 VPWR VGND sg13g2_decap_8
Xhold9 _040_ VPWR VGND net22 sg13g2_dlygate4sd3_1
X_069_ genblk1\[1\].csa.hsum2 _033_ _035_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_16 VPWR VGND sg13g2_fill_1
X_085_ net41 net18 _047_ VPWR VGND sg13g2_xor2_1
XFILLER_0_84 VPWR VGND sg13g2_decap_8
X_068_ net34 VPWR _001_ VGND _033_ _034_ sg13g2_o21ai_1
Xfanout1 net2 net1 VPWR VGND sg13g2_buf_8
X_084_ net18 genblk1\[4\].csa.y _046_ VPWR VGND sg13g2_nor2_1
XFILLER_0_30 VPWR VGND sg13g2_decap_8
X_067_ net40 net33 _035_ VPWR VGND sg13g2_xor2_1
Xfanout2 net3 net2 VPWR VGND sg13g2_buf_8
X_119_ _013_ VGND VPWR genblk1\[1\].csa.hsum2 csa0.y clknet_2_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_12_94 VPWR VGND sg13g2_decap_8
X_083_ _045_ net12 net8 VPWR VGND sg13g2_nand2_1
X_118_ _012_ VGND VPWR _008_ tcmp.z clknet_2_2__leaf_clk sg13g2_dfrbpq_1
X_066_ net33 genblk1\[1\].csa.y _034_ VPWR VGND sg13g2_nor2_1
XFILLER_3_106 VPWR VGND sg13g2_fill_1
XFILLER_7_4 VPWR VGND sg13g2_fill_1
X_082_ _044_ net18 genblk1\[4\].csa.y VPWR VGND sg13g2_nand2_1
X_065_ _033_ net12 net5 VPWR VGND sg13g2_nand2_1
XFILLER_0_98 VPWR VGND sg13g2_decap_8
X_117_ _011_ VGND VPWR _007_ genblk1\[6\].csa.y clknet_2_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_12_74 VPWR VGND sg13g2_decap_4
XFILLER_12_52 VPWR VGND sg13g2_fill_1
X_081_ genblk1\[3\].csa.hsum2 _041_ _043_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_53 VPWR VGND sg13g2_decap_8
X_064_ _032_ net33 genblk1\[1\].csa.y VPWR VGND sg13g2_nand2_1
X_116_ _010_ VGND VPWR net17 csa0.sc clknet_2_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_3_11 VPWR VGND sg13g2_fill_2
XFILLER_12_42 VPWR VGND sg13g2_fill_1
X_080_ net22 VPWR _003_ VGND _041_ _042_ sg13g2_o21ai_1
X_063_ _007_ net14 _031_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_23 VPWR VGND sg13g2_decap_8
X_115_ _009_ VGND VPWR csa0.hsum2 net13 clknet_2_1__leaf_clk sg13g2_dfrbpq_1
.ends

