VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spm
  CLASS BLOCK ;
  FOREIGN spm ;
  ORIGIN 0.000 0.000 ;
  SIZE 62.920 BY 81.640 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal1 ;
        RECT 24.460 14.490 26.660 64.480 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 5.540 33.820 57.340 36.020 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TopMetal1 ;
        RECT 18.260 14.900 20.460 64.890 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 5.540 27.620 57.340 29.820 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal3 ;
        RECT 62.520 21.220 62.920 21.620 ;
    END
  END clk
  PIN p
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 62.520 37.180 62.920 37.580 ;
    END
  END p
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.340 0.400 57.740 ;
    END
  END rst
  PIN x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 62.520 31.300 62.920 31.700 ;
    END
  END x[0]
  PIN x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 34.840 0.000 35.240 0.400 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 28.780 0.400 29.180 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 34.660 0.400 35.060 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 62.520 43.900 62.920 44.300 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 35.800 81.240 36.200 81.640 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 20.440 81.240 20.840 81.640 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 45.580 0.400 45.980 ;
    END
  END x[7]
  PIN y
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.500 0.400 56.900 ;
    END
  END y
  OBS
      LAYER GatPoly ;
        RECT 5.760 14.970 57.120 64.410 ;
      LAYER Metal1 ;
        RECT 5.760 14.900 57.120 64.480 ;
      LAYER Metal2 ;
        RECT 5.655 81.030 20.230 81.240 ;
        RECT 21.050 81.030 35.590 81.240 ;
        RECT 36.410 81.030 57.225 81.240 ;
        RECT 5.655 0.610 57.225 81.030 ;
        RECT 5.655 0.400 34.630 0.610 ;
        RECT 35.450 0.400 57.225 0.610 ;
      LAYER Metal3 ;
        RECT 0.400 57.950 62.520 69.400 ;
        RECT 0.610 57.130 62.520 57.950 ;
        RECT 0.400 57.110 62.520 57.130 ;
        RECT 0.610 56.290 62.520 57.110 ;
        RECT 0.400 46.190 62.520 56.290 ;
        RECT 0.610 45.370 62.520 46.190 ;
        RECT 0.400 44.510 62.520 45.370 ;
        RECT 0.400 43.690 62.310 44.510 ;
        RECT 0.400 37.790 62.520 43.690 ;
        RECT 0.400 36.970 62.310 37.790 ;
        RECT 0.400 35.270 62.520 36.970 ;
        RECT 0.610 34.450 62.520 35.270 ;
        RECT 0.400 31.910 62.520 34.450 ;
        RECT 0.400 31.090 62.310 31.910 ;
        RECT 0.400 29.390 62.520 31.090 ;
        RECT 0.610 28.570 62.520 29.390 ;
        RECT 0.400 21.830 62.520 28.570 ;
        RECT 0.400 21.010 62.310 21.830 ;
        RECT 0.400 6.200 62.520 21.010 ;
      LAYER Metal4 ;
        RECT 9.495 14.975 31.785 64.405 ;
      LAYER Metal5 ;
        RECT 9.455 14.810 31.825 64.570 ;
  END
END spm
END LIBRARY

